-- 500 variable assigns in 2 processes. GHC works here.

entity main is
end entity main;

architecture arch of main is
	signal clk : integer := 0;
	constant CYCLES : integer := 1000;
begin

	main: process(clk)
--{{{
		variable a0502 : integer;
		variable a0503 : integer;
		variable a0504 : integer;
		variable a0505 : integer;
		variable a0506 : integer;
		variable a0507 : integer;
		variable a0508 : integer;
		variable a0509 : integer;
		variable a0510 : integer;
		variable a0511 : integer;
		variable a0512 : integer;
		variable a0513 : integer;
		variable a0514 : integer;
		variable a0515 : integer;
		variable a0516 : integer;
		variable a0517 : integer;
		variable a0518 : integer;
		variable a0519 : integer;
		variable a0520 : integer;
		variable a0521 : integer;
		variable a0522 : integer;
		variable a0523 : integer;
		variable a0524 : integer;
		variable a0525 : integer;
		variable a0526 : integer;
		variable a0527 : integer;
		variable a0528 : integer;
		variable a0529 : integer;
		variable a0530 : integer;
		variable a0531 : integer;
		variable a0532 : integer;
		variable a0533 : integer;
		variable a0534 : integer;
		variable a0535 : integer;
		variable a0536 : integer;
		variable a0537 : integer;
		variable a0538 : integer;
		variable a0539 : integer;
		variable a0540 : integer;
		variable a0541 : integer;
		variable a0542 : integer;
		variable a0543 : integer;
		variable a0544 : integer;
		variable a0545 : integer;
		variable a0546 : integer;
		variable a0547 : integer;
		variable a0548 : integer;
		variable a0549 : integer;
		variable a0550 : integer;
		variable a0551 : integer;
		variable a0552 : integer;
		variable a0553 : integer;
		variable a0554 : integer;
		variable a0555 : integer;
		variable a0556 : integer;
		variable a0557 : integer;
		variable a0558 : integer;
		variable a0559 : integer;
		variable a0560 : integer;
		variable a0561 : integer;
		variable a0562 : integer;
		variable a0563 : integer;
		variable a0564 : integer;
		variable a0565 : integer;
		variable a0566 : integer;
		variable a0567 : integer;
		variable a0568 : integer;
		variable a0569 : integer;
		variable a0570 : integer;
		variable a0571 : integer;
		variable a0572 : integer;
		variable a0573 : integer;
		variable a0574 : integer;
		variable a0575 : integer;
		variable a0576 : integer;
		variable a0577 : integer;
		variable a0578 : integer;
		variable a0579 : integer;
		variable a0580 : integer;
		variable a0581 : integer;
		variable a0582 : integer;
		variable a0583 : integer;
		variable a0584 : integer;
		variable a0585 : integer;
		variable a0586 : integer;
		variable a0587 : integer;
		variable a0588 : integer;
		variable a0589 : integer;
		variable a0590 : integer;
		variable a0591 : integer;
		variable a0592 : integer;
		variable a0593 : integer;
		variable a0594 : integer;
		variable a0595 : integer;
		variable a0596 : integer;
		variable a0597 : integer;
		variable a0598 : integer;
		variable a0599 : integer;
		variable a0600 : integer;
		variable a0601 : integer;
		variable a0602 : integer;
		variable a0603 : integer;
		variable a0604 : integer;
		variable a0605 : integer;
		variable a0606 : integer;
		variable a0607 : integer;
		variable a0608 : integer;
		variable a0609 : integer;
		variable a0610 : integer;
		variable a0611 : integer;
		variable a0612 : integer;
		variable a0613 : integer;
		variable a0614 : integer;
		variable a0615 : integer;
		variable a0616 : integer;
		variable a0617 : integer;
		variable a0618 : integer;
		variable a0619 : integer;
		variable a0620 : integer;
		variable a0621 : integer;
		variable a0622 : integer;
		variable a0623 : integer;
		variable a0624 : integer;
		variable a0625 : integer;
		variable a0626 : integer;
		variable a0627 : integer;
		variable a0628 : integer;
		variable a0629 : integer;
		variable a0630 : integer;
		variable a0631 : integer;
		variable a0632 : integer;
		variable a0633 : integer;
		variable a0634 : integer;
		variable a0635 : integer;
		variable a0636 : integer;
		variable a0637 : integer;
		variable a0638 : integer;
		variable a0639 : integer;
		variable a0640 : integer;
		variable a0641 : integer;
		variable a0642 : integer;
		variable a0643 : integer;
		variable a0644 : integer;
		variable a0645 : integer;
		variable a0646 : integer;
		variable a0647 : integer;
		variable a0648 : integer;
		variable a0649 : integer;
		variable a0650 : integer;
		variable a0651 : integer;
		variable a0652 : integer;
		variable a0653 : integer;
		variable a0654 : integer;
		variable a0655 : integer;
		variable a0656 : integer;
		variable a0657 : integer;
		variable a0658 : integer;
		variable a0659 : integer;
		variable a0660 : integer;
		variable a0661 : integer;
		variable a0662 : integer;
		variable a0663 : integer;
		variable a0664 : integer;
		variable a0665 : integer;
		variable a0666 : integer;
		variable a0667 : integer;
		variable a0668 : integer;
		variable a0669 : integer;
		variable a0670 : integer;
		variable a0671 : integer;
		variable a0672 : integer;
		variable a0673 : integer;
		variable a0674 : integer;
		variable a0675 : integer;
		variable a0676 : integer;
		variable a0677 : integer;
		variable a0678 : integer;
		variable a0679 : integer;
		variable a0680 : integer;
		variable a0681 : integer;
		variable a0682 : integer;
		variable a0683 : integer;
		variable a0684 : integer;
		variable a0685 : integer;
		variable a0686 : integer;
		variable a0687 : integer;
		variable a0688 : integer;
		variable a0689 : integer;
		variable a0690 : integer;
		variable a0691 : integer;
		variable a0692 : integer;
		variable a0693 : integer;
		variable a0694 : integer;
		variable a0695 : integer;
		variable a0696 : integer;
		variable a0697 : integer;
		variable a0698 : integer;
		variable a0699 : integer;
		variable a0700 : integer;
		variable a0701 : integer;
		variable a0702 : integer;
		variable a0703 : integer;
		variable a0704 : integer;
		variable a0705 : integer;
		variable a0706 : integer;
		variable a0707 : integer;
		variable a0708 : integer;
		variable a0709 : integer;
		variable a0710 : integer;
		variable a0711 : integer;
		variable a0712 : integer;
		variable a0713 : integer;
		variable a0714 : integer;
		variable a0715 : integer;
		variable a0716 : integer;
		variable a0717 : integer;
		variable a0718 : integer;
		variable a0719 : integer;
		variable a0720 : integer;
		variable a0721 : integer;
		variable a0722 : integer;
		variable a0723 : integer;
		variable a0724 : integer;
		variable a0725 : integer;
		variable a0726 : integer;
		variable a0727 : integer;
		variable a0728 : integer;
		variable a0729 : integer;
		variable a0730 : integer;
		variable a0731 : integer;
		variable a0732 : integer;
		variable a0733 : integer;
		variable a0734 : integer;
		variable a0735 : integer;
		variable a0736 : integer;
		variable a0737 : integer;
		variable a0738 : integer;
		variable a0739 : integer;
		variable a0740 : integer;
		variable a0741 : integer;
		variable a0742 : integer;
		variable a0743 : integer;
		variable a0744 : integer;
		variable a0745 : integer;
		variable a0746 : integer;
		variable a0747 : integer;
		variable a0748 : integer;
		variable a0749 : integer;
		variable a0750 : integer;
		variable a0751 : integer;
		variable a0752 : integer;
		variable a0753 : integer;
		variable a0754 : integer;
		variable a0755 : integer;
		variable a0756 : integer;
		variable a0757 : integer;
		variable a0758 : integer;
		variable a0759 : integer;
		variable a0760 : integer;
		variable a0761 : integer;
		variable a0762 : integer;
		variable a0763 : integer;
		variable a0764 : integer;
		variable a0765 : integer;
		variable a0766 : integer;
		variable a0767 : integer;
		variable a0768 : integer;
		variable a0769 : integer;
		variable a0770 : integer;
		variable a0771 : integer;
		variable a0772 : integer;
		variable a0773 : integer;
		variable a0774 : integer;
		variable a0775 : integer;
		variable a0776 : integer;
		variable a0777 : integer;
		variable a0778 : integer;
		variable a0779 : integer;
		variable a0780 : integer;
		variable a0781 : integer;
		variable a0782 : integer;
		variable a0783 : integer;
		variable a0784 : integer;
		variable a0785 : integer;
		variable a0786 : integer;
		variable a0787 : integer;
		variable a0788 : integer;
		variable a0789 : integer;
		variable a0790 : integer;
		variable a0791 : integer;
		variable a0792 : integer;
		variable a0793 : integer;
		variable a0794 : integer;
		variable a0795 : integer;
		variable a0796 : integer;
		variable a0797 : integer;
		variable a0798 : integer;
		variable a0799 : integer;
		variable a0800 : integer;
		variable a0801 : integer;
		variable a0802 : integer;
		variable a0803 : integer;
		variable a0804 : integer;
		variable a0805 : integer;
		variable a0806 : integer;
		variable a0807 : integer;
		variable a0808 : integer;
		variable a0809 : integer;
		variable a0810 : integer;
		variable a0811 : integer;
		variable a0812 : integer;
		variable a0813 : integer;
		variable a0814 : integer;
		variable a0815 : integer;
		variable a0816 : integer;
		variable a0817 : integer;
		variable a0818 : integer;
		variable a0819 : integer;
		variable a0820 : integer;
		variable a0821 : integer;
		variable a0822 : integer;
		variable a0823 : integer;
		variable a0824 : integer;
		variable a0825 : integer;
		variable a0826 : integer;
		variable a0827 : integer;
		variable a0828 : integer;
		variable a0829 : integer;
		variable a0830 : integer;
		variable a0831 : integer;
		variable a0832 : integer;
		variable a0833 : integer;
		variable a0834 : integer;
		variable a0835 : integer;
		variable a0836 : integer;
		variable a0837 : integer;
		variable a0838 : integer;
		variable a0839 : integer;
		variable a0840 : integer;
		variable a0841 : integer;
		variable a0842 : integer;
		variable a0843 : integer;
		variable a0844 : integer;
		variable a0845 : integer;
		variable a0846 : integer;
		variable a0847 : integer;
		variable a0848 : integer;
		variable a0849 : integer;
		variable a0850 : integer;
		variable a0851 : integer;
		variable a0852 : integer;
		variable a0853 : integer;
		variable a0854 : integer;
		variable a0855 : integer;
		variable a0856 : integer;
		variable a0857 : integer;
		variable a0858 : integer;
		variable a0859 : integer;
		variable a0860 : integer;
		variable a0861 : integer;
		variable a0862 : integer;
		variable a0863 : integer;
		variable a0864 : integer;
		variable a0865 : integer;
		variable a0866 : integer;
		variable a0867 : integer;
		variable a0868 : integer;
		variable a0869 : integer;
		variable a0870 : integer;
		variable a0871 : integer;
		variable a0872 : integer;
		variable a0873 : integer;
		variable a0874 : integer;
		variable a0875 : integer;
		variable a0876 : integer;
		variable a0877 : integer;
		variable a0878 : integer;
		variable a0879 : integer;
		variable a0880 : integer;
		variable a0881 : integer;
		variable a0882 : integer;
		variable a0883 : integer;
		variable a0884 : integer;
		variable a0885 : integer;
		variable a0886 : integer;
		variable a0887 : integer;
		variable a0888 : integer;
		variable a0889 : integer;
		variable a0890 : integer;
		variable a0891 : integer;
		variable a0892 : integer;
		variable a0893 : integer;
		variable a0894 : integer;
		variable a0895 : integer;
		variable a0896 : integer;
		variable a0897 : integer;
		variable a0898 : integer;
		variable a0899 : integer;
		variable a0900 : integer;
		variable a0901 : integer;
		variable a0902 : integer;
		variable a0903 : integer;
		variable a0904 : integer;
		variable a0905 : integer;
		variable a0906 : integer;
		variable a0907 : integer;
		variable a0908 : integer;
		variable a0909 : integer;
		variable a0910 : integer;
		variable a0911 : integer;
		variable a0912 : integer;
		variable a0913 : integer;
		variable a0914 : integer;
		variable a0915 : integer;
		variable a0916 : integer;
		variable a0917 : integer;
		variable a0918 : integer;
		variable a0919 : integer;
		variable a0920 : integer;
		variable a0921 : integer;
		variable a0922 : integer;
		variable a0923 : integer;
		variable a0924 : integer;
		variable a0925 : integer;
		variable a0926 : integer;
		variable a0927 : integer;
		variable a0928 : integer;
		variable a0929 : integer;
		variable a0930 : integer;
		variable a0931 : integer;
		variable a0932 : integer;
		variable a0933 : integer;
		variable a0934 : integer;
		variable a0935 : integer;
		variable a0936 : integer;
		variable a0937 : integer;
		variable a0938 : integer;
		variable a0939 : integer;
		variable a0940 : integer;
		variable a0941 : integer;
		variable a0942 : integer;
		variable a0943 : integer;
		variable a0944 : integer;
		variable a0945 : integer;
		variable a0946 : integer;
		variable a0947 : integer;
		variable a0948 : integer;
		variable a0949 : integer;
		variable a0950 : integer;
		variable a0951 : integer;
		variable a0952 : integer;
		variable a0953 : integer;
		variable a0954 : integer;
		variable a0955 : integer;
		variable a0956 : integer;
		variable a0957 : integer;
		variable a0958 : integer;
		variable a0959 : integer;
		variable a0960 : integer;
		variable a0961 : integer;
		variable a0962 : integer;
		variable a0963 : integer;
		variable a0964 : integer;
		variable a0965 : integer;
		variable a0966 : integer;
		variable a0967 : integer;
		variable a0968 : integer;
		variable a0969 : integer;
		variable a0970 : integer;
		variable a0971 : integer;
		variable a0972 : integer;
		variable a0973 : integer;
		variable a0974 : integer;
		variable a0975 : integer;
		variable a0976 : integer;
		variable a0977 : integer;
		variable a0978 : integer;
		variable a0979 : integer;
		variable a0980 : integer;
		variable a0981 : integer;
		variable a0982 : integer;
		variable a0983 : integer;
		variable a0984 : integer;
		variable a0985 : integer;
		variable a0986 : integer;
		variable a0987 : integer;
		variable a0988 : integer;
		variable a0989 : integer;
		variable a0990 : integer;
		variable a0991 : integer;
		variable a0992 : integer;
		variable a0993 : integer;
		variable a0994 : integer;
		variable a0995 : integer;
		variable a0996 : integer;
		variable a0997 : integer;
		variable a0998 : integer;
		variable a0999 : integer;
		variable a1000 : integer;
	begin
		a0502 := 502;
		a0503 := 503;
		a0504 := 504;
		a0505 := 505;
		a0506 := 506;
		a0507 := 507;
		a0508 := 508;
		a0509 := 509;
		a0510 := 510;
		a0511 := 511;
		a0512 := 512;
		a0513 := 513;
		a0514 := 514;
		a0515 := 515;
		a0516 := 516;
		a0517 := 517;
		a0518 := 518;
		a0519 := 519;
		a0520 := 520;
		a0521 := 521;
		a0522 := 522;
		a0523 := 523;
		a0524 := 524;
		a0525 := 525;
		a0526 := 526;
		a0527 := 527;
		a0528 := 528;
		a0529 := 529;
		a0530 := 530;
		a0531 := 531;
		a0532 := 532;
		a0533 := 533;
		a0534 := 534;
		a0535 := 535;
		a0536 := 536;
		a0537 := 537;
		a0538 := 538;
		a0539 := 539;
		a0540 := 540;
		a0541 := 541;
		a0542 := 542;
		a0543 := 543;
		a0544 := 544;
		a0545 := 545;
		a0546 := 546;
		a0547 := 547;
		a0548 := 548;
		a0549 := 549;
		a0550 := 550;
		a0551 := 551;
		a0552 := 552;
		a0553 := 553;
		a0554 := 554;
		a0555 := 555;
		a0556 := 556;
		a0557 := 557;
		a0558 := 558;
		a0559 := 559;
		a0560 := 560;
		a0561 := 561;
		a0562 := 562;
		a0563 := 563;
		a0564 := 564;
		a0565 := 565;
		a0566 := 566;
		a0567 := 567;
		a0568 := 568;
		a0569 := 569;
		a0570 := 570;
		a0571 := 571;
		a0572 := 572;
		a0573 := 573;
		a0574 := 574;
		a0575 := 575;
		a0576 := 576;
		a0577 := 577;
		a0578 := 578;
		a0579 := 579;
		a0580 := 580;
		a0581 := 581;
		a0582 := 582;
		a0583 := 583;
		a0584 := 584;
		a0585 := 585;
		a0586 := 586;
		a0587 := 587;
		a0588 := 588;
		a0589 := 589;
		a0590 := 590;
		a0591 := 591;
		a0592 := 592;
		a0593 := 593;
		a0594 := 594;
		a0595 := 595;
		a0596 := 596;
		a0597 := 597;
		a0598 := 598;
		a0599 := 599;
		a0600 := 600;
		a0601 := 601;
		a0602 := 602;
		a0603 := 603;
		a0604 := 604;
		a0605 := 605;
		a0606 := 606;
		a0607 := 607;
		a0608 := 608;
		a0609 := 609;
		a0610 := 610;
		a0611 := 611;
		a0612 := 612;
		a0613 := 613;
		a0614 := 614;
		a0615 := 615;
		a0616 := 616;
		a0617 := 617;
		a0618 := 618;
		a0619 := 619;
		a0620 := 620;
		a0621 := 621;
		a0622 := 622;
		a0623 := 623;
		a0624 := 624;
		a0625 := 625;
		a0626 := 626;
		a0627 := 627;
		a0628 := 628;
		a0629 := 629;
		a0630 := 630;
		a0631 := 631;
		a0632 := 632;
		a0633 := 633;
		a0634 := 634;
		a0635 := 635;
		a0636 := 636;
		a0637 := 637;
		a0638 := 638;
		a0639 := 639;
		a0640 := 640;
		a0641 := 641;
		a0642 := 642;
		a0643 := 643;
		a0644 := 644;
		a0645 := 645;
		a0646 := 646;
		a0647 := 647;
		a0648 := 648;
		a0649 := 649;
		a0650 := 650;
		a0651 := 651;
		a0652 := 652;
		a0653 := 653;
		a0654 := 654;
		a0655 := 655;
		a0656 := 656;
		a0657 := 657;
		a0658 := 658;
		a0659 := 659;
		a0660 := 660;
		a0661 := 661;
		a0662 := 662;
		a0663 := 663;
		a0664 := 664;
		a0665 := 665;
		a0666 := 666;
		a0667 := 667;
		a0668 := 668;
		a0669 := 669;
		a0670 := 670;
		a0671 := 671;
		a0672 := 672;
		a0673 := 673;
		a0674 := 674;
		a0675 := 675;
		a0676 := 676;
		a0677 := 677;
		a0678 := 678;
		a0679 := 679;
		a0680 := 680;
		a0681 := 681;
		a0682 := 682;
		a0683 := 683;
		a0684 := 684;
		a0685 := 685;
		a0686 := 686;
		a0687 := 687;
		a0688 := 688;
		a0689 := 689;
		a0690 := 690;
		a0691 := 691;
		a0692 := 692;
		a0693 := 693;
		a0694 := 694;
		a0695 := 695;
		a0696 := 696;
		a0697 := 697;
		a0698 := 698;
		a0699 := 699;
		a0700 := 700;
		a0701 := 701;
		a0702 := 702;
		a0703 := 703;
		a0704 := 704;
		a0705 := 705;
		a0706 := 706;
		a0707 := 707;
		a0708 := 708;
		a0709 := 709;
		a0710 := 710;
		a0711 := 711;
		a0712 := 712;
		a0713 := 713;
		a0714 := 714;
		a0715 := 715;
		a0716 := 716;
		a0717 := 717;
		a0718 := 718;
		a0719 := 719;
		a0720 := 720;
		a0721 := 721;
		a0722 := 722;
		a0723 := 723;
		a0724 := 724;
		a0725 := 725;
		a0726 := 726;
		a0727 := 727;
		a0728 := 728;
		a0729 := 729;
		a0730 := 730;
		a0731 := 731;
		a0732 := 732;
		a0733 := 733;
		a0734 := 734;
		a0735 := 735;
		a0736 := 736;
		a0737 := 737;
		a0738 := 738;
		a0739 := 739;
		a0740 := 740;
		a0741 := 741;
		a0742 := 742;
		a0743 := 743;
		a0744 := 744;
		a0745 := 745;
		a0746 := 746;
		a0747 := 747;
		a0748 := 748;
		a0749 := 749;
		a0750 := 750;
		a0751 := 751;
		a0752 := 752;
		a0753 := 753;
		a0754 := 754;
		a0755 := 755;
		a0756 := 756;
		a0757 := 757;
		a0758 := 758;
		a0759 := 759;
		a0760 := 760;
		a0761 := 761;
		a0762 := 762;
		a0763 := 763;
		a0764 := 764;
		a0765 := 765;
		a0766 := 766;
		a0767 := 767;
		a0768 := 768;
		a0769 := 769;
		a0770 := 770;
		a0771 := 771;
		a0772 := 772;
		a0773 := 773;
		a0774 := 774;
		a0775 := 775;
		a0776 := 776;
		a0777 := 777;
		a0778 := 778;
		a0779 := 779;
		a0780 := 780;
		a0781 := 781;
		a0782 := 782;
		a0783 := 783;
		a0784 := 784;
		a0785 := 785;
		a0786 := 786;
		a0787 := 787;
		a0788 := 788;
		a0789 := 789;
		a0790 := 790;
		a0791 := 791;
		a0792 := 792;
		a0793 := 793;
		a0794 := 794;
		a0795 := 795;
		a0796 := 796;
		a0797 := 797;
		a0798 := 798;
		a0799 := 799;
		a0800 := 800;
		a0801 := 801;
		a0802 := 802;
		a0803 := 803;
		a0804 := 804;
		a0805 := 805;
		a0806 := 806;
		a0807 := 807;
		a0808 := 808;
		a0809 := 809;
		a0810 := 810;
		a0811 := 811;
		a0812 := 812;
		a0813 := 813;
		a0814 := 814;
		a0815 := 815;
		a0816 := 816;
		a0817 := 817;
		a0818 := 818;
		a0819 := 819;
		a0820 := 820;
		a0821 := 821;
		a0822 := 822;
		a0823 := 823;
		a0824 := 824;
		a0825 := 825;
		a0826 := 826;
		a0827 := 827;
		a0828 := 828;
		a0829 := 829;
		a0830 := 830;
		a0831 := 831;
		a0832 := 832;
		a0833 := 833;
		a0834 := 834;
		a0835 := 835;
		a0836 := 836;
		a0837 := 837;
		a0838 := 838;
		a0839 := 839;
		a0840 := 840;
		a0841 := 841;
		a0842 := 842;
		a0843 := 843;
		a0844 := 844;
		a0845 := 845;
		a0846 := 846;
		a0847 := 847;
		a0848 := 848;
		a0849 := 849;
		a0850 := 850;
		a0851 := 851;
		a0852 := 852;
		a0853 := 853;
		a0854 := 854;
		a0855 := 855;
		a0856 := 856;
		a0857 := 857;
		a0858 := 858;
		a0859 := 859;
		a0860 := 860;
		a0861 := 861;
		a0862 := 862;
		a0863 := 863;
		a0864 := 864;
		a0865 := 865;
		a0866 := 866;
		a0867 := 867;
		a0868 := 868;
		a0869 := 869;
		a0870 := 870;
		a0871 := 871;
		a0872 := 872;
		a0873 := 873;
		a0874 := 874;
		a0875 := 875;
		a0876 := 876;
		a0877 := 877;
		a0878 := 878;
		a0879 := 879;
		a0880 := 880;
		a0881 := 881;
		a0882 := 882;
		a0883 := 883;
		a0884 := 884;
		a0885 := 885;
		a0886 := 886;
		a0887 := 887;
		a0888 := 888;
		a0889 := 889;
		a0890 := 890;
		a0891 := 891;
		a0892 := 892;
		a0893 := 893;
		a0894 := 894;
		a0895 := 895;
		a0896 := 896;
		a0897 := 897;
		a0898 := 898;
		a0899 := 899;
		a0900 := 900;
		a0901 := 901;
		a0902 := 902;
		a0903 := 903;
		a0904 := 904;
		a0905 := 905;
		a0906 := 906;
		a0907 := 907;
		a0908 := 908;
		a0909 := 909;
		a0910 := 910;
		a0911 := 911;
		a0912 := 912;
		a0913 := 913;
		a0914 := 914;
		a0915 := 915;
		a0916 := 916;
		a0917 := 917;
		a0918 := 918;
		a0919 := 919;
		a0920 := 920;
		a0921 := 921;
		a0922 := 922;
		a0923 := 923;
		a0924 := 924;
		a0925 := 925;
		a0926 := 926;
		a0927 := 927;
		a0928 := 928;
		a0929 := 929;
		a0930 := 930;
		a0931 := 931;
		a0932 := 932;
		a0933 := 933;
		a0934 := 934;
		a0935 := 935;
		a0936 := 936;
		a0937 := 937;
		a0938 := 938;
		a0939 := 939;
		a0940 := 940;
		a0941 := 941;
		a0942 := 942;
		a0943 := 943;
		a0944 := 944;
		a0945 := 945;
		a0946 := 946;
		a0947 := 947;
		a0948 := 948;
		a0949 := 949;
		a0950 := 950;
		a0951 := 951;
		a0952 := 952;
		a0953 := 953;
		a0954 := 954;
		a0955 := 955;
		a0956 := 956;
		a0957 := 957;
		a0958 := 958;
		a0959 := 959;
		a0960 := 960;
		a0961 := 961;
		a0962 := 962;
		a0963 := 963;
		a0964 := 964;
		a0965 := 965;
		a0966 := 966;
		a0967 := 967;
		a0968 := 968;
		a0969 := 969;
		a0970 := 970;
		a0971 := 971;
		a0972 := 972;
		a0973 := 973;
		a0974 := 974;
		a0975 := 975;
		a0976 := 976;
		a0977 := 977;
		a0978 := 978;
		a0979 := 979;
		a0980 := 980;
		a0981 := 981;
		a0982 := 982;
		a0983 := 983;
		a0984 := 984;
		a0985 := 985;
		a0986 := 986;
		a0987 := 987;
		a0988 := 988;
		a0989 := 989;
		a0990 := 990;
		a0991 := 991;
		a0992 := 992;
		a0993 := 993;
		a0994 := 994;
		a0995 := 995;
		a0996 := 996;
		a0997 := 997;
		a0998 := 998;
		a0999 := 999;
		a1000 := 1000;
        -- report "tick";
--}}}
    end process;

	main2: process(clk)
--{{{
		variable a0502 : integer;
		variable a0503 : integer;
		variable a0504 : integer;
		variable a0505 : integer;
		variable a0506 : integer;
		variable a0507 : integer;
		variable a0508 : integer;
		variable a0509 : integer;
		variable a0510 : integer;
		variable a0511 : integer;
		variable a0512 : integer;
		variable a0513 : integer;
		variable a0514 : integer;
		variable a0515 : integer;
		variable a0516 : integer;
		variable a0517 : integer;
		variable a0518 : integer;
		variable a0519 : integer;
		variable a0520 : integer;
		variable a0521 : integer;
		variable a0522 : integer;
		variable a0523 : integer;
		variable a0524 : integer;
		variable a0525 : integer;
		variable a0526 : integer;
		variable a0527 : integer;
		variable a0528 : integer;
		variable a0529 : integer;
		variable a0530 : integer;
		variable a0531 : integer;
		variable a0532 : integer;
		variable a0533 : integer;
		variable a0534 : integer;
		variable a0535 : integer;
		variable a0536 : integer;
		variable a0537 : integer;
		variable a0538 : integer;
		variable a0539 : integer;
		variable a0540 : integer;
		variable a0541 : integer;
		variable a0542 : integer;
		variable a0543 : integer;
		variable a0544 : integer;
		variable a0545 : integer;
		variable a0546 : integer;
		variable a0547 : integer;
		variable a0548 : integer;
		variable a0549 : integer;
		variable a0550 : integer;
		variable a0551 : integer;
		variable a0552 : integer;
		variable a0553 : integer;
		variable a0554 : integer;
		variable a0555 : integer;
		variable a0556 : integer;
		variable a0557 : integer;
		variable a0558 : integer;
		variable a0559 : integer;
		variable a0560 : integer;
		variable a0561 : integer;
		variable a0562 : integer;
		variable a0563 : integer;
		variable a0564 : integer;
		variable a0565 : integer;
		variable a0566 : integer;
		variable a0567 : integer;
		variable a0568 : integer;
		variable a0569 : integer;
		variable a0570 : integer;
		variable a0571 : integer;
		variable a0572 : integer;
		variable a0573 : integer;
		variable a0574 : integer;
		variable a0575 : integer;
		variable a0576 : integer;
		variable a0577 : integer;
		variable a0578 : integer;
		variable a0579 : integer;
		variable a0580 : integer;
		variable a0581 : integer;
		variable a0582 : integer;
		variable a0583 : integer;
		variable a0584 : integer;
		variable a0585 : integer;
		variable a0586 : integer;
		variable a0587 : integer;
		variable a0588 : integer;
		variable a0589 : integer;
		variable a0590 : integer;
		variable a0591 : integer;
		variable a0592 : integer;
		variable a0593 : integer;
		variable a0594 : integer;
		variable a0595 : integer;
		variable a0596 : integer;
		variable a0597 : integer;
		variable a0598 : integer;
		variable a0599 : integer;
		variable a0600 : integer;
		variable a0601 : integer;
		variable a0602 : integer;
		variable a0603 : integer;
		variable a0604 : integer;
		variable a0605 : integer;
		variable a0606 : integer;
		variable a0607 : integer;
		variable a0608 : integer;
		variable a0609 : integer;
		variable a0610 : integer;
		variable a0611 : integer;
		variable a0612 : integer;
		variable a0613 : integer;
		variable a0614 : integer;
		variable a0615 : integer;
		variable a0616 : integer;
		variable a0617 : integer;
		variable a0618 : integer;
		variable a0619 : integer;
		variable a0620 : integer;
		variable a0621 : integer;
		variable a0622 : integer;
		variable a0623 : integer;
		variable a0624 : integer;
		variable a0625 : integer;
		variable a0626 : integer;
		variable a0627 : integer;
		variable a0628 : integer;
		variable a0629 : integer;
		variable a0630 : integer;
		variable a0631 : integer;
		variable a0632 : integer;
		variable a0633 : integer;
		variable a0634 : integer;
		variable a0635 : integer;
		variable a0636 : integer;
		variable a0637 : integer;
		variable a0638 : integer;
		variable a0639 : integer;
		variable a0640 : integer;
		variable a0641 : integer;
		variable a0642 : integer;
		variable a0643 : integer;
		variable a0644 : integer;
		variable a0645 : integer;
		variable a0646 : integer;
		variable a0647 : integer;
		variable a0648 : integer;
		variable a0649 : integer;
		variable a0650 : integer;
		variable a0651 : integer;
		variable a0652 : integer;
		variable a0653 : integer;
		variable a0654 : integer;
		variable a0655 : integer;
		variable a0656 : integer;
		variable a0657 : integer;
		variable a0658 : integer;
		variable a0659 : integer;
		variable a0660 : integer;
		variable a0661 : integer;
		variable a0662 : integer;
		variable a0663 : integer;
		variable a0664 : integer;
		variable a0665 : integer;
		variable a0666 : integer;
		variable a0667 : integer;
		variable a0668 : integer;
		variable a0669 : integer;
		variable a0670 : integer;
		variable a0671 : integer;
		variable a0672 : integer;
		variable a0673 : integer;
		variable a0674 : integer;
		variable a0675 : integer;
		variable a0676 : integer;
		variable a0677 : integer;
		variable a0678 : integer;
		variable a0679 : integer;
		variable a0680 : integer;
		variable a0681 : integer;
		variable a0682 : integer;
		variable a0683 : integer;
		variable a0684 : integer;
		variable a0685 : integer;
		variable a0686 : integer;
		variable a0687 : integer;
		variable a0688 : integer;
		variable a0689 : integer;
		variable a0690 : integer;
		variable a0691 : integer;
		variable a0692 : integer;
		variable a0693 : integer;
		variable a0694 : integer;
		variable a0695 : integer;
		variable a0696 : integer;
		variable a0697 : integer;
		variable a0698 : integer;
		variable a0699 : integer;
		variable a0700 : integer;
		variable a0701 : integer;
		variable a0702 : integer;
		variable a0703 : integer;
		variable a0704 : integer;
		variable a0705 : integer;
		variable a0706 : integer;
		variable a0707 : integer;
		variable a0708 : integer;
		variable a0709 : integer;
		variable a0710 : integer;
		variable a0711 : integer;
		variable a0712 : integer;
		variable a0713 : integer;
		variable a0714 : integer;
		variable a0715 : integer;
		variable a0716 : integer;
		variable a0717 : integer;
		variable a0718 : integer;
		variable a0719 : integer;
		variable a0720 : integer;
		variable a0721 : integer;
		variable a0722 : integer;
		variable a0723 : integer;
		variable a0724 : integer;
		variable a0725 : integer;
		variable a0726 : integer;
		variable a0727 : integer;
		variable a0728 : integer;
		variable a0729 : integer;
		variable a0730 : integer;
		variable a0731 : integer;
		variable a0732 : integer;
		variable a0733 : integer;
		variable a0734 : integer;
		variable a0735 : integer;
		variable a0736 : integer;
		variable a0737 : integer;
		variable a0738 : integer;
		variable a0739 : integer;
		variable a0740 : integer;
		variable a0741 : integer;
		variable a0742 : integer;
		variable a0743 : integer;
		variable a0744 : integer;
		variable a0745 : integer;
		variable a0746 : integer;
		variable a0747 : integer;
		variable a0748 : integer;
		variable a0749 : integer;
		variable a0750 : integer;
		variable a0751 : integer;
		variable a0752 : integer;
		variable a0753 : integer;
		variable a0754 : integer;
		variable a0755 : integer;
		variable a0756 : integer;
		variable a0757 : integer;
		variable a0758 : integer;
		variable a0759 : integer;
		variable a0760 : integer;
		variable a0761 : integer;
		variable a0762 : integer;
		variable a0763 : integer;
		variable a0764 : integer;
		variable a0765 : integer;
		variable a0766 : integer;
		variable a0767 : integer;
		variable a0768 : integer;
		variable a0769 : integer;
		variable a0770 : integer;
		variable a0771 : integer;
		variable a0772 : integer;
		variable a0773 : integer;
		variable a0774 : integer;
		variable a0775 : integer;
		variable a0776 : integer;
		variable a0777 : integer;
		variable a0778 : integer;
		variable a0779 : integer;
		variable a0780 : integer;
		variable a0781 : integer;
		variable a0782 : integer;
		variable a0783 : integer;
		variable a0784 : integer;
		variable a0785 : integer;
		variable a0786 : integer;
		variable a0787 : integer;
		variable a0788 : integer;
		variable a0789 : integer;
		variable a0790 : integer;
		variable a0791 : integer;
		variable a0792 : integer;
		variable a0793 : integer;
		variable a0794 : integer;
		variable a0795 : integer;
		variable a0796 : integer;
		variable a0797 : integer;
		variable a0798 : integer;
		variable a0799 : integer;
		variable a0800 : integer;
		variable a0801 : integer;
		variable a0802 : integer;
		variable a0803 : integer;
		variable a0804 : integer;
		variable a0805 : integer;
		variable a0806 : integer;
		variable a0807 : integer;
		variable a0808 : integer;
		variable a0809 : integer;
		variable a0810 : integer;
		variable a0811 : integer;
		variable a0812 : integer;
		variable a0813 : integer;
		variable a0814 : integer;
		variable a0815 : integer;
		variable a0816 : integer;
		variable a0817 : integer;
		variable a0818 : integer;
		variable a0819 : integer;
		variable a0820 : integer;
		variable a0821 : integer;
		variable a0822 : integer;
		variable a0823 : integer;
		variable a0824 : integer;
		variable a0825 : integer;
		variable a0826 : integer;
		variable a0827 : integer;
		variable a0828 : integer;
		variable a0829 : integer;
		variable a0830 : integer;
		variable a0831 : integer;
		variable a0832 : integer;
		variable a0833 : integer;
		variable a0834 : integer;
		variable a0835 : integer;
		variable a0836 : integer;
		variable a0837 : integer;
		variable a0838 : integer;
		variable a0839 : integer;
		variable a0840 : integer;
		variable a0841 : integer;
		variable a0842 : integer;
		variable a0843 : integer;
		variable a0844 : integer;
		variable a0845 : integer;
		variable a0846 : integer;
		variable a0847 : integer;
		variable a0848 : integer;
		variable a0849 : integer;
		variable a0850 : integer;
		variable a0851 : integer;
		variable a0852 : integer;
		variable a0853 : integer;
		variable a0854 : integer;
		variable a0855 : integer;
		variable a0856 : integer;
		variable a0857 : integer;
		variable a0858 : integer;
		variable a0859 : integer;
		variable a0860 : integer;
		variable a0861 : integer;
		variable a0862 : integer;
		variable a0863 : integer;
		variable a0864 : integer;
		variable a0865 : integer;
		variable a0866 : integer;
		variable a0867 : integer;
		variable a0868 : integer;
		variable a0869 : integer;
		variable a0870 : integer;
		variable a0871 : integer;
		variable a0872 : integer;
		variable a0873 : integer;
		variable a0874 : integer;
		variable a0875 : integer;
		variable a0876 : integer;
		variable a0877 : integer;
		variable a0878 : integer;
		variable a0879 : integer;
		variable a0880 : integer;
		variable a0881 : integer;
		variable a0882 : integer;
		variable a0883 : integer;
		variable a0884 : integer;
		variable a0885 : integer;
		variable a0886 : integer;
		variable a0887 : integer;
		variable a0888 : integer;
		variable a0889 : integer;
		variable a0890 : integer;
		variable a0891 : integer;
		variable a0892 : integer;
		variable a0893 : integer;
		variable a0894 : integer;
		variable a0895 : integer;
		variable a0896 : integer;
		variable a0897 : integer;
		variable a0898 : integer;
		variable a0899 : integer;
		variable a0900 : integer;
		variable a0901 : integer;
		variable a0902 : integer;
		variable a0903 : integer;
		variable a0904 : integer;
		variable a0905 : integer;
		variable a0906 : integer;
		variable a0907 : integer;
		variable a0908 : integer;
		variable a0909 : integer;
		variable a0910 : integer;
		variable a0911 : integer;
		variable a0912 : integer;
		variable a0913 : integer;
		variable a0914 : integer;
		variable a0915 : integer;
		variable a0916 : integer;
		variable a0917 : integer;
		variable a0918 : integer;
		variable a0919 : integer;
		variable a0920 : integer;
		variable a0921 : integer;
		variable a0922 : integer;
		variable a0923 : integer;
		variable a0924 : integer;
		variable a0925 : integer;
		variable a0926 : integer;
		variable a0927 : integer;
		variable a0928 : integer;
		variable a0929 : integer;
		variable a0930 : integer;
		variable a0931 : integer;
		variable a0932 : integer;
		variable a0933 : integer;
		variable a0934 : integer;
		variable a0935 : integer;
		variable a0936 : integer;
		variable a0937 : integer;
		variable a0938 : integer;
		variable a0939 : integer;
		variable a0940 : integer;
		variable a0941 : integer;
		variable a0942 : integer;
		variable a0943 : integer;
		variable a0944 : integer;
		variable a0945 : integer;
		variable a0946 : integer;
		variable a0947 : integer;
		variable a0948 : integer;
		variable a0949 : integer;
		variable a0950 : integer;
		variable a0951 : integer;
		variable a0952 : integer;
		variable a0953 : integer;
		variable a0954 : integer;
		variable a0955 : integer;
		variable a0956 : integer;
		variable a0957 : integer;
		variable a0958 : integer;
		variable a0959 : integer;
		variable a0960 : integer;
		variable a0961 : integer;
		variable a0962 : integer;
		variable a0963 : integer;
		variable a0964 : integer;
		variable a0965 : integer;
		variable a0966 : integer;
		variable a0967 : integer;
		variable a0968 : integer;
		variable a0969 : integer;
		variable a0970 : integer;
		variable a0971 : integer;
		variable a0972 : integer;
		variable a0973 : integer;
		variable a0974 : integer;
		variable a0975 : integer;
		variable a0976 : integer;
		variable a0977 : integer;
		variable a0978 : integer;
		variable a0979 : integer;
		variable a0980 : integer;
		variable a0981 : integer;
		variable a0982 : integer;
		variable a0983 : integer;
		variable a0984 : integer;
		variable a0985 : integer;
		variable a0986 : integer;
		variable a0987 : integer;
		variable a0988 : integer;
		variable a0989 : integer;
		variable a0990 : integer;
		variable a0991 : integer;
		variable a0992 : integer;
		variable a0993 : integer;
		variable a0994 : integer;
		variable a0995 : integer;
		variable a0996 : integer;
		variable a0997 : integer;
		variable a0998 : integer;
		variable a0999 : integer;
		variable a1000 : integer;
	begin
		a0502 := 502;
		a0503 := 503;
		a0504 := 504;
		a0505 := 505;
		a0506 := 506;
		a0507 := 507;
		a0508 := 508;
		a0509 := 509;
		a0510 := 510;
		a0511 := 511;
		a0512 := 512;
		a0513 := 513;
		a0514 := 514;
		a0515 := 515;
		a0516 := 516;
		a0517 := 517;
		a0518 := 518;
		a0519 := 519;
		a0520 := 520;
		a0521 := 521;
		a0522 := 522;
		a0523 := 523;
		a0524 := 524;
		a0525 := 525;
		a0526 := 526;
		a0527 := 527;
		a0528 := 528;
		a0529 := 529;
		a0530 := 530;
		a0531 := 531;
		a0532 := 532;
		a0533 := 533;
		a0534 := 534;
		a0535 := 535;
		a0536 := 536;
		a0537 := 537;
		a0538 := 538;
		a0539 := 539;
		a0540 := 540;
		a0541 := 541;
		a0542 := 542;
		a0543 := 543;
		a0544 := 544;
		a0545 := 545;
		a0546 := 546;
		a0547 := 547;
		a0548 := 548;
		a0549 := 549;
		a0550 := 550;
		a0551 := 551;
		a0552 := 552;
		a0553 := 553;
		a0554 := 554;
		a0555 := 555;
		a0556 := 556;
		a0557 := 557;
		a0558 := 558;
		a0559 := 559;
		a0560 := 560;
		a0561 := 561;
		a0562 := 562;
		a0563 := 563;
		a0564 := 564;
		a0565 := 565;
		a0566 := 566;
		a0567 := 567;
		a0568 := 568;
		a0569 := 569;
		a0570 := 570;
		a0571 := 571;
		a0572 := 572;
		a0573 := 573;
		a0574 := 574;
		a0575 := 575;
		a0576 := 576;
		a0577 := 577;
		a0578 := 578;
		a0579 := 579;
		a0580 := 580;
		a0581 := 581;
		a0582 := 582;
		a0583 := 583;
		a0584 := 584;
		a0585 := 585;
		a0586 := 586;
		a0587 := 587;
		a0588 := 588;
		a0589 := 589;
		a0590 := 590;
		a0591 := 591;
		a0592 := 592;
		a0593 := 593;
		a0594 := 594;
		a0595 := 595;
		a0596 := 596;
		a0597 := 597;
		a0598 := 598;
		a0599 := 599;
		a0600 := 600;
		a0601 := 601;
		a0602 := 602;
		a0603 := 603;
		a0604 := 604;
		a0605 := 605;
		a0606 := 606;
		a0607 := 607;
		a0608 := 608;
		a0609 := 609;
		a0610 := 610;
		a0611 := 611;
		a0612 := 612;
		a0613 := 613;
		a0614 := 614;
		a0615 := 615;
		a0616 := 616;
		a0617 := 617;
		a0618 := 618;
		a0619 := 619;
		a0620 := 620;
		a0621 := 621;
		a0622 := 622;
		a0623 := 623;
		a0624 := 624;
		a0625 := 625;
		a0626 := 626;
		a0627 := 627;
		a0628 := 628;
		a0629 := 629;
		a0630 := 630;
		a0631 := 631;
		a0632 := 632;
		a0633 := 633;
		a0634 := 634;
		a0635 := 635;
		a0636 := 636;
		a0637 := 637;
		a0638 := 638;
		a0639 := 639;
		a0640 := 640;
		a0641 := 641;
		a0642 := 642;
		a0643 := 643;
		a0644 := 644;
		a0645 := 645;
		a0646 := 646;
		a0647 := 647;
		a0648 := 648;
		a0649 := 649;
		a0650 := 650;
		a0651 := 651;
		a0652 := 652;
		a0653 := 653;
		a0654 := 654;
		a0655 := 655;
		a0656 := 656;
		a0657 := 657;
		a0658 := 658;
		a0659 := 659;
		a0660 := 660;
		a0661 := 661;
		a0662 := 662;
		a0663 := 663;
		a0664 := 664;
		a0665 := 665;
		a0666 := 666;
		a0667 := 667;
		a0668 := 668;
		a0669 := 669;
		a0670 := 670;
		a0671 := 671;
		a0672 := 672;
		a0673 := 673;
		a0674 := 674;
		a0675 := 675;
		a0676 := 676;
		a0677 := 677;
		a0678 := 678;
		a0679 := 679;
		a0680 := 680;
		a0681 := 681;
		a0682 := 682;
		a0683 := 683;
		a0684 := 684;
		a0685 := 685;
		a0686 := 686;
		a0687 := 687;
		a0688 := 688;
		a0689 := 689;
		a0690 := 690;
		a0691 := 691;
		a0692 := 692;
		a0693 := 693;
		a0694 := 694;
		a0695 := 695;
		a0696 := 696;
		a0697 := 697;
		a0698 := 698;
		a0699 := 699;
		a0700 := 700;
		a0701 := 701;
		a0702 := 702;
		a0703 := 703;
		a0704 := 704;
		a0705 := 705;
		a0706 := 706;
		a0707 := 707;
		a0708 := 708;
		a0709 := 709;
		a0710 := 710;
		a0711 := 711;
		a0712 := 712;
		a0713 := 713;
		a0714 := 714;
		a0715 := 715;
		a0716 := 716;
		a0717 := 717;
		a0718 := 718;
		a0719 := 719;
		a0720 := 720;
		a0721 := 721;
		a0722 := 722;
		a0723 := 723;
		a0724 := 724;
		a0725 := 725;
		a0726 := 726;
		a0727 := 727;
		a0728 := 728;
		a0729 := 729;
		a0730 := 730;
		a0731 := 731;
		a0732 := 732;
		a0733 := 733;
		a0734 := 734;
		a0735 := 735;
		a0736 := 736;
		a0737 := 737;
		a0738 := 738;
		a0739 := 739;
		a0740 := 740;
		a0741 := 741;
		a0742 := 742;
		a0743 := 743;
		a0744 := 744;
		a0745 := 745;
		a0746 := 746;
		a0747 := 747;
		a0748 := 748;
		a0749 := 749;
		a0750 := 750;
		a0751 := 751;
		a0752 := 752;
		a0753 := 753;
		a0754 := 754;
		a0755 := 755;
		a0756 := 756;
		a0757 := 757;
		a0758 := 758;
		a0759 := 759;
		a0760 := 760;
		a0761 := 761;
		a0762 := 762;
		a0763 := 763;
		a0764 := 764;
		a0765 := 765;
		a0766 := 766;
		a0767 := 767;
		a0768 := 768;
		a0769 := 769;
		a0770 := 770;
		a0771 := 771;
		a0772 := 772;
		a0773 := 773;
		a0774 := 774;
		a0775 := 775;
		a0776 := 776;
		a0777 := 777;
		a0778 := 778;
		a0779 := 779;
		a0780 := 780;
		a0781 := 781;
		a0782 := 782;
		a0783 := 783;
		a0784 := 784;
		a0785 := 785;
		a0786 := 786;
		a0787 := 787;
		a0788 := 788;
		a0789 := 789;
		a0790 := 790;
		a0791 := 791;
		a0792 := 792;
		a0793 := 793;
		a0794 := 794;
		a0795 := 795;
		a0796 := 796;
		a0797 := 797;
		a0798 := 798;
		a0799 := 799;
		a0800 := 800;
		a0801 := 801;
		a0802 := 802;
		a0803 := 803;
		a0804 := 804;
		a0805 := 805;
		a0806 := 806;
		a0807 := 807;
		a0808 := 808;
		a0809 := 809;
		a0810 := 810;
		a0811 := 811;
		a0812 := 812;
		a0813 := 813;
		a0814 := 814;
		a0815 := 815;
		a0816 := 816;
		a0817 := 817;
		a0818 := 818;
		a0819 := 819;
		a0820 := 820;
		a0821 := 821;
		a0822 := 822;
		a0823 := 823;
		a0824 := 824;
		a0825 := 825;
		a0826 := 826;
		a0827 := 827;
		a0828 := 828;
		a0829 := 829;
		a0830 := 830;
		a0831 := 831;
		a0832 := 832;
		a0833 := 833;
		a0834 := 834;
		a0835 := 835;
		a0836 := 836;
		a0837 := 837;
		a0838 := 838;
		a0839 := 839;
		a0840 := 840;
		a0841 := 841;
		a0842 := 842;
		a0843 := 843;
		a0844 := 844;
		a0845 := 845;
		a0846 := 846;
		a0847 := 847;
		a0848 := 848;
		a0849 := 849;
		a0850 := 850;
		a0851 := 851;
		a0852 := 852;
		a0853 := 853;
		a0854 := 854;
		a0855 := 855;
		a0856 := 856;
		a0857 := 857;
		a0858 := 858;
		a0859 := 859;
		a0860 := 860;
		a0861 := 861;
		a0862 := 862;
		a0863 := 863;
		a0864 := 864;
		a0865 := 865;
		a0866 := 866;
		a0867 := 867;
		a0868 := 868;
		a0869 := 869;
		a0870 := 870;
		a0871 := 871;
		a0872 := 872;
		a0873 := 873;
		a0874 := 874;
		a0875 := 875;
		a0876 := 876;
		a0877 := 877;
		a0878 := 878;
		a0879 := 879;
		a0880 := 880;
		a0881 := 881;
		a0882 := 882;
		a0883 := 883;
		a0884 := 884;
		a0885 := 885;
		a0886 := 886;
		a0887 := 887;
		a0888 := 888;
		a0889 := 889;
		a0890 := 890;
		a0891 := 891;
		a0892 := 892;
		a0893 := 893;
		a0894 := 894;
		a0895 := 895;
		a0896 := 896;
		a0897 := 897;
		a0898 := 898;
		a0899 := 899;
		a0900 := 900;
		a0901 := 901;
		a0902 := 902;
		a0903 := 903;
		a0904 := 904;
		a0905 := 905;
		a0906 := 906;
		a0907 := 907;
		a0908 := 908;
		a0909 := 909;
		a0910 := 910;
		a0911 := 911;
		a0912 := 912;
		a0913 := 913;
		a0914 := 914;
		a0915 := 915;
		a0916 := 916;
		a0917 := 917;
		a0918 := 918;
		a0919 := 919;
		a0920 := 920;
		a0921 := 921;
		a0922 := 922;
		a0923 := 923;
		a0924 := 924;
		a0925 := 925;
		a0926 := 926;
		a0927 := 927;
		a0928 := 928;
		a0929 := 929;
		a0930 := 930;
		a0931 := 931;
		a0932 := 932;
		a0933 := 933;
		a0934 := 934;
		a0935 := 935;
		a0936 := 936;
		a0937 := 937;
		a0938 := 938;
		a0939 := 939;
		a0940 := 940;
		a0941 := 941;
		a0942 := 942;
		a0943 := 943;
		a0944 := 944;
		a0945 := 945;
		a0946 := 946;
		a0947 := 947;
		a0948 := 948;
		a0949 := 949;
		a0950 := 950;
		a0951 := 951;
		a0952 := 952;
		a0953 := 953;
		a0954 := 954;
		a0955 := 955;
		a0956 := 956;
		a0957 := 957;
		a0958 := 958;
		a0959 := 959;
		a0960 := 960;
		a0961 := 961;
		a0962 := 962;
		a0963 := 963;
		a0964 := 964;
		a0965 := 965;
		a0966 := 966;
		a0967 := 967;
		a0968 := 968;
		a0969 := 969;
		a0970 := 970;
		a0971 := 971;
		a0972 := 972;
		a0973 := 973;
		a0974 := 974;
		a0975 := 975;
		a0976 := 976;
		a0977 := 977;
		a0978 := 978;
		a0979 := 979;
		a0980 := 980;
		a0981 := 981;
		a0982 := 982;
		a0983 := 983;
		a0984 := 984;
		a0985 := 985;
		a0986 := 986;
		a0987 := 987;
		a0988 := 988;
		a0989 := 989;
		a0990 := 990;
		a0991 := 991;
		a0992 := 992;
		a0993 := 993;
		a0994 := 994;
		a0995 := 995;
		a0996 := 996;
		a0997 := 997;
		a0998 := 998;
		a0999 := 999;
		a1000 := 1000;
        -- report "tick";
--}}}
    end process;

	terminator : process(clk)
	begin
		if clk >= CYCLES then
			assert false report "end of simulation" severity failure;
		-- else
		-- 	report "tick";
		end if;
	end process;

	clk <= (clk+1) after 1 us;
end;
