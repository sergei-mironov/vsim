entity ENT00001_Test_Bench is
end entity ENT00001_Test_Bench;

architecture arch of ENT00001_Test_Bench is
	signal clk : integer := 0;
	constant CYCLES : integer := 10000;
	-- {{{
	signal a0001 : integer;
	signal a0002 : integer;
	signal a0003 : integer;
	signal a0004 : integer;
	signal a0005 : integer;
	signal a0006 : integer;
	signal a0007 : integer;
	signal a0008 : integer;
	signal a0009 : integer;
	signal a0010 : integer;
	signal a0011 : integer;
	signal a0012 : integer;
	signal a0013 : integer;
	signal a0014 : integer;
	signal a0015 : integer;
	signal a0016 : integer;
	signal a0017 : integer;
	signal a0018 : integer;
	signal a0019 : integer;
	signal a0020 : integer;
	signal a0021 : integer;
	signal a0022 : integer;
	signal a0023 : integer;
	signal a0024 : integer;
	signal a0025 : integer;
	signal a0026 : integer;
	signal a0027 : integer;
	signal a0028 : integer;
	signal a0029 : integer;
	signal a0030 : integer;
	signal a0031 : integer;
	signal a0032 : integer;
	signal a0033 : integer;
	signal a0034 : integer;
	signal a0035 : integer;
	signal a0036 : integer;
	signal a0037 : integer;
	signal a0038 : integer;
	signal a0039 : integer;
	signal a0040 : integer;
	signal a0041 : integer;
	signal a0042 : integer;
	signal a0043 : integer;
	signal a0044 : integer;
	signal a0045 : integer;
	signal a0046 : integer;
	signal a0047 : integer;
	signal a0048 : integer;
	signal a0049 : integer;
	signal a0050 : integer;
	signal a0051 : integer;
	signal a0052 : integer;
	signal a0053 : integer;
	signal a0054 : integer;
	signal a0055 : integer;
	signal a0056 : integer;
	signal a0057 : integer;
	signal a0058 : integer;
	signal a0059 : integer;
	signal a0060 : integer;
	signal a0061 : integer;
	signal a0062 : integer;
	signal a0063 : integer;
	signal a0064 : integer;
	signal a0065 : integer;
	signal a0066 : integer;
	signal a0067 : integer;
	signal a0068 : integer;
	signal a0069 : integer;
	signal a0070 : integer;
	signal a0071 : integer;
	signal a0072 : integer;
	signal a0073 : integer;
	signal a0074 : integer;
	signal a0075 : integer;
	signal a0076 : integer;
	signal a0077 : integer;
	signal a0078 : integer;
	signal a0079 : integer;
	signal a0080 : integer;
	signal a0081 : integer;
	signal a0082 : integer;
	signal a0083 : integer;
	signal a0084 : integer;
	signal a0085 : integer;
	signal a0086 : integer;
	signal a0087 : integer;
	signal a0088 : integer;
	signal a0089 : integer;
	signal a0090 : integer;
	signal a0091 : integer;
	signal a0092 : integer;
	signal a0093 : integer;
	signal a0094 : integer;
	signal a0095 : integer;
	signal a0096 : integer;
	signal a0097 : integer;
	signal a0098 : integer;
	signal a0099 : integer;
	signal a0100 : integer;
	signal a0101 : integer;
	signal a0102 : integer;
	signal a0103 : integer;
	signal a0104 : integer;
	signal a0105 : integer;
	signal a0106 : integer;
	signal a0107 : integer;
	signal a0108 : integer;
	signal a0109 : integer;
	signal a0110 : integer;
	signal a0111 : integer;
	signal a0112 : integer;
	signal a0113 : integer;
	signal a0114 : integer;
	signal a0115 : integer;
	signal a0116 : integer;
	signal a0117 : integer;
	signal a0118 : integer;
	signal a0119 : integer;
	signal a0120 : integer;
	signal a0121 : integer;
	signal a0122 : integer;
	signal a0123 : integer;
	signal a0124 : integer;
	signal a0125 : integer;
	signal a0126 : integer;
	signal a0127 : integer;
	signal a0128 : integer;
	signal a0129 : integer;
	signal a0130 : integer;
	signal a0131 : integer;
	signal a0132 : integer;
	signal a0133 : integer;
	signal a0134 : integer;
	signal a0135 : integer;
	signal a0136 : integer;
	signal a0137 : integer;
	signal a0138 : integer;
	signal a0139 : integer;
	signal a0140 : integer;
	signal a0141 : integer;
	signal a0142 : integer;
	signal a0143 : integer;
	signal a0144 : integer;
	signal a0145 : integer;
	signal a0146 : integer;
	signal a0147 : integer;
	signal a0148 : integer;
	signal a0149 : integer;
	signal a0150 : integer;
	signal a0151 : integer;
	signal a0152 : integer;
	signal a0153 : integer;
	signal a0154 : integer;
	signal a0155 : integer;
	signal a0156 : integer;
	signal a0157 : integer;
	signal a0158 : integer;
	signal a0159 : integer;
	signal a0160 : integer;
	signal a0161 : integer;
	signal a0162 : integer;
	signal a0163 : integer;
	signal a0164 : integer;
	signal a0165 : integer;
	signal a0166 : integer;
	signal a0167 : integer;
	signal a0168 : integer;
	signal a0169 : integer;
	signal a0170 : integer;
	signal a0171 : integer;
	signal a0172 : integer;
	signal a0173 : integer;
	signal a0174 : integer;
	signal a0175 : integer;
	signal a0176 : integer;
	signal a0177 : integer;
	signal a0178 : integer;
	signal a0179 : integer;
	signal a0180 : integer;
	signal a0181 : integer;
	signal a0182 : integer;
	signal a0183 : integer;
	signal a0184 : integer;
	signal a0185 : integer;
	signal a0186 : integer;
	signal a0187 : integer;
	signal a0188 : integer;
	signal a0189 : integer;
	signal a0190 : integer;
	signal a0191 : integer;
	signal a0192 : integer;
	signal a0193 : integer;
	signal a0194 : integer;
	signal a0195 : integer;
	signal a0196 : integer;
	signal a0197 : integer;
	signal a0198 : integer;
	signal a0199 : integer;
	signal a0200 : integer;
	signal a0201 : integer;
	signal a0202 : integer;
	signal a0203 : integer;
	signal a0204 : integer;
	signal a0205 : integer;
	signal a0206 : integer;
	signal a0207 : integer;
	signal a0208 : integer;
	signal a0209 : integer;
	signal a0210 : integer;
	signal a0211 : integer;
	signal a0212 : integer;
	signal a0213 : integer;
	signal a0214 : integer;
	signal a0215 : integer;
	signal a0216 : integer;
	signal a0217 : integer;
	signal a0218 : integer;
	signal a0219 : integer;
	signal a0220 : integer;
	signal a0221 : integer;
	signal a0222 : integer;
	signal a0223 : integer;
	signal a0224 : integer;
	signal a0225 : integer;
	signal a0226 : integer;
	signal a0227 : integer;
	signal a0228 : integer;
	signal a0229 : integer;
	signal a0230 : integer;
	signal a0231 : integer;
	signal a0232 : integer;
	signal a0233 : integer;
	signal a0234 : integer;
	signal a0235 : integer;
	signal a0236 : integer;
	signal a0237 : integer;
	signal a0238 : integer;
	signal a0239 : integer;
	signal a0240 : integer;
	signal a0241 : integer;
	signal a0242 : integer;
	signal a0243 : integer;
	signal a0244 : integer;
	signal a0245 : integer;
	signal a0246 : integer;
	signal a0247 : integer;
	signal a0248 : integer;
	signal a0249 : integer;
	signal a0250 : integer;
	signal a0251 : integer;
	signal a0252 : integer;
	signal a0253 : integer;
	signal a0254 : integer;
	signal a0255 : integer;
	signal a0256 : integer;
	signal a0257 : integer;
	signal a0258 : integer;
	signal a0259 : integer;
	signal a0260 : integer;
	signal a0261 : integer;
	signal a0262 : integer;
	signal a0263 : integer;
	signal a0264 : integer;
	signal a0265 : integer;
	signal a0266 : integer;
	signal a0267 : integer;
	signal a0268 : integer;
	signal a0269 : integer;
	signal a0270 : integer;
	signal a0271 : integer;
	signal a0272 : integer;
	signal a0273 : integer;
	signal a0274 : integer;
	signal a0275 : integer;
	signal a0276 : integer;
	signal a0277 : integer;
	signal a0278 : integer;
	signal a0279 : integer;
	signal a0280 : integer;
	signal a0281 : integer;
	signal a0282 : integer;
	signal a0283 : integer;
	signal a0284 : integer;
	signal a0285 : integer;
	signal a0286 : integer;
	signal a0287 : integer;
	signal a0288 : integer;
	signal a0289 : integer;
	signal a0290 : integer;
	signal a0291 : integer;
	signal a0292 : integer;
	signal a0293 : integer;
	signal a0294 : integer;
	signal a0295 : integer;
	signal a0296 : integer;
	signal a0297 : integer;
	signal a0298 : integer;
	signal a0299 : integer;
	signal a0300 : integer;
	signal a0301 : integer;
	signal a0302 : integer;
	signal a0303 : integer;
	signal a0304 : integer;
	signal a0305 : integer;
	signal a0306 : integer;
	signal a0307 : integer;
	signal a0308 : integer;
	signal a0309 : integer;
	signal a0310 : integer;
	signal a0311 : integer;
	signal a0312 : integer;
	signal a0313 : integer;
	signal a0314 : integer;
	signal a0315 : integer;
	signal a0316 : integer;
	signal a0317 : integer;
	signal a0318 : integer;
	signal a0319 : integer;
	signal a0320 : integer;
	signal a0321 : integer;
	signal a0322 : integer;
	signal a0323 : integer;
	signal a0324 : integer;
	signal a0325 : integer;
	signal a0326 : integer;
	signal a0327 : integer;
	signal a0328 : integer;
	signal a0329 : integer;
	signal a0330 : integer;
	signal a0331 : integer;
	signal a0332 : integer;
	signal a0333 : integer;
	signal a0334 : integer;
	signal a0335 : integer;
	signal a0336 : integer;
	signal a0337 : integer;
	signal a0338 : integer;
	signal a0339 : integer;
	signal a0340 : integer;
	signal a0341 : integer;
	signal a0342 : integer;
	signal a0343 : integer;
	signal a0344 : integer;
	signal a0345 : integer;
	signal a0346 : integer;
	signal a0347 : integer;
	signal a0348 : integer;
	signal a0349 : integer;
	signal a0350 : integer;
	signal a0351 : integer;
	signal a0352 : integer;
	signal a0353 : integer;
	signal a0354 : integer;
	signal a0355 : integer;
	signal a0356 : integer;
	signal a0357 : integer;
	signal a0358 : integer;
	signal a0359 : integer;
	signal a0360 : integer;
	signal a0361 : integer;
	signal a0362 : integer;
	signal a0363 : integer;
	signal a0364 : integer;
	signal a0365 : integer;
	signal a0366 : integer;
	signal a0367 : integer;
	signal a0368 : integer;
	signal a0369 : integer;
	signal a0370 : integer;
	signal a0371 : integer;
	signal a0372 : integer;
	signal a0373 : integer;
	signal a0374 : integer;
	signal a0375 : integer;
	signal a0376 : integer;
	signal a0377 : integer;
	signal a0378 : integer;
	signal a0379 : integer;
	signal a0380 : integer;
	signal a0381 : integer;
	signal a0382 : integer;
	signal a0383 : integer;
	signal a0384 : integer;
	signal a0385 : integer;
	signal a0386 : integer;
	signal a0387 : integer;
	signal a0388 : integer;
	signal a0389 : integer;
	signal a0390 : integer;
	signal a0391 : integer;
	signal a0392 : integer;
	signal a0393 : integer;
	signal a0394 : integer;
	signal a0395 : integer;
	signal a0396 : integer;
	signal a0397 : integer;
	signal a0398 : integer;
	signal a0399 : integer;
	signal a0400 : integer;
	signal a0401 : integer;
	signal a0402 : integer;
	signal a0403 : integer;
	signal a0404 : integer;
	signal a0405 : integer;
	signal a0406 : integer;
	signal a0407 : integer;
	signal a0408 : integer;
	signal a0409 : integer;
	signal a0410 : integer;
	signal a0411 : integer;
	signal a0412 : integer;
	signal a0413 : integer;
	signal a0414 : integer;
	signal a0415 : integer;
	signal a0416 : integer;
	signal a0417 : integer;
	signal a0418 : integer;
	signal a0419 : integer;
	signal a0420 : integer;
	signal a0421 : integer;
	signal a0422 : integer;
	signal a0423 : integer;
	signal a0424 : integer;
	signal a0425 : integer;
	signal a0426 : integer;
	signal a0427 : integer;
	signal a0428 : integer;
	signal a0429 : integer;
	signal a0430 : integer;
	signal a0431 : integer;
	signal a0432 : integer;
	signal a0433 : integer;
	signal a0434 : integer;
	signal a0435 : integer;
	signal a0436 : integer;
	signal a0437 : integer;
	signal a0438 : integer;
	signal a0439 : integer;
	signal a0440 : integer;
	signal a0441 : integer;
	signal a0442 : integer;
	signal a0443 : integer;
	signal a0444 : integer;
	signal a0445 : integer;
	signal a0446 : integer;
	signal a0447 : integer;
	signal a0448 : integer;
	signal a0449 : integer;
	signal a0450 : integer;
	signal a0451 : integer;
	signal a0452 : integer;
	signal a0453 : integer;
	signal a0454 : integer;
	signal a0455 : integer;
	signal a0456 : integer;
	signal a0457 : integer;
	signal a0458 : integer;
	signal a0459 : integer;
	signal a0460 : integer;
	signal a0461 : integer;
	signal a0462 : integer;
	signal a0463 : integer;
	signal a0464 : integer;
	signal a0465 : integer;
	signal a0466 : integer;
	signal a0467 : integer;
	signal a0468 : integer;
	signal a0469 : integer;
	signal a0470 : integer;
	signal a0471 : integer;
	signal a0472 : integer;
	signal a0473 : integer;
	signal a0474 : integer;
	signal a0475 : integer;
	signal a0476 : integer;
	signal a0477 : integer;
	signal a0478 : integer;
	signal a0479 : integer;
	signal a0480 : integer;
	signal a0481 : integer;
	signal a0482 : integer;
	signal a0483 : integer;
	signal a0484 : integer;
	signal a0485 : integer;
	signal a0486 : integer;
	signal a0487 : integer;
	signal a0488 : integer;
	signal a0489 : integer;
	signal a0490 : integer;
	signal a0491 : integer;
	signal a0492 : integer;
	signal a0493 : integer;
	signal a0494 : integer;
	signal a0495 : integer;
	signal a0496 : integer;
	signal a0497 : integer;
	signal a0498 : integer;
	signal a0499 : integer;
	signal a0500 : integer;
	signal a0501 : integer;
	signal a0502 : integer;
	signal a0503 : integer;
	signal a0504 : integer;
	signal a0505 : integer;
	signal a0506 : integer;
	signal a0507 : integer;
	signal a0508 : integer;
	signal a0509 : integer;
	signal a0510 : integer;
	signal a0511 : integer;
	signal a0512 : integer;
	signal a0513 : integer;
	signal a0514 : integer;
	signal a0515 : integer;
	signal a0516 : integer;
	signal a0517 : integer;
	signal a0518 : integer;
	signal a0519 : integer;
	signal a0520 : integer;
	signal a0521 : integer;
	signal a0522 : integer;
	signal a0523 : integer;
	signal a0524 : integer;
	signal a0525 : integer;
	signal a0526 : integer;
	signal a0527 : integer;
	signal a0528 : integer;
	signal a0529 : integer;
	signal a0530 : integer;
	signal a0531 : integer;
	signal a0532 : integer;
	signal a0533 : integer;
	signal a0534 : integer;
	signal a0535 : integer;
	signal a0536 : integer;
	signal a0537 : integer;
	signal a0538 : integer;
	signal a0539 : integer;
	signal a0540 : integer;
	signal a0541 : integer;
	signal a0542 : integer;
	signal a0543 : integer;
	signal a0544 : integer;
	signal a0545 : integer;
	signal a0546 : integer;
	signal a0547 : integer;
	signal a0548 : integer;
	signal a0549 : integer;
	signal a0550 : integer;
	signal a0551 : integer;
	signal a0552 : integer;
	signal a0553 : integer;
	signal a0554 : integer;
	signal a0555 : integer;
	signal a0556 : integer;
	signal a0557 : integer;
	signal a0558 : integer;
	signal a0559 : integer;
	signal a0560 : integer;
	signal a0561 : integer;
	signal a0562 : integer;
	signal a0563 : integer;
	signal a0564 : integer;
	signal a0565 : integer;
	signal a0566 : integer;
	signal a0567 : integer;
	signal a0568 : integer;
	signal a0569 : integer;
	signal a0570 : integer;
	signal a0571 : integer;
	signal a0572 : integer;
	signal a0573 : integer;
	signal a0574 : integer;
	signal a0575 : integer;
	signal a0576 : integer;
	signal a0577 : integer;
	signal a0578 : integer;
	signal a0579 : integer;
	signal a0580 : integer;
	signal a0581 : integer;
	signal a0582 : integer;
	signal a0583 : integer;
	signal a0584 : integer;
	signal a0585 : integer;
	signal a0586 : integer;
	signal a0587 : integer;
	signal a0588 : integer;
	signal a0589 : integer;
	signal a0590 : integer;
	signal a0591 : integer;
	signal a0592 : integer;
	signal a0593 : integer;
	signal a0594 : integer;
	signal a0595 : integer;
	signal a0596 : integer;
	signal a0597 : integer;
	signal a0598 : integer;
	signal a0599 : integer;
	signal a0600 : integer;
	signal a0601 : integer;
	signal a0602 : integer;
	signal a0603 : integer;
	signal a0604 : integer;
	signal a0605 : integer;
	signal a0606 : integer;
	signal a0607 : integer;
	signal a0608 : integer;
	signal a0609 : integer;
	signal a0610 : integer;
	signal a0611 : integer;
	signal a0612 : integer;
	signal a0613 : integer;
	signal a0614 : integer;
	signal a0615 : integer;
	signal a0616 : integer;
	signal a0617 : integer;
	signal a0618 : integer;
	signal a0619 : integer;
	signal a0620 : integer;
	signal a0621 : integer;
	signal a0622 : integer;
	signal a0623 : integer;
	signal a0624 : integer;
	signal a0625 : integer;
	signal a0626 : integer;
	signal a0627 : integer;
	signal a0628 : integer;
	signal a0629 : integer;
	signal a0630 : integer;
	signal a0631 : integer;
	signal a0632 : integer;
	signal a0633 : integer;
	signal a0634 : integer;
	signal a0635 : integer;
	signal a0636 : integer;
	signal a0637 : integer;
	signal a0638 : integer;
	signal a0639 : integer;
	signal a0640 : integer;
	signal a0641 : integer;
	signal a0642 : integer;
	signal a0643 : integer;
	signal a0644 : integer;
	signal a0645 : integer;
	signal a0646 : integer;
	signal a0647 : integer;
	signal a0648 : integer;
	signal a0649 : integer;
	signal a0650 : integer;
	signal a0651 : integer;
	signal a0652 : integer;
	signal a0653 : integer;
	signal a0654 : integer;
	signal a0655 : integer;
	signal a0656 : integer;
	signal a0657 : integer;
	signal a0658 : integer;
	signal a0659 : integer;
	signal a0660 : integer;
	signal a0661 : integer;
	signal a0662 : integer;
	signal a0663 : integer;
	signal a0664 : integer;
	signal a0665 : integer;
	signal a0666 : integer;
	signal a0667 : integer;
	signal a0668 : integer;
	signal a0669 : integer;
	signal a0670 : integer;
	signal a0671 : integer;
	signal a0672 : integer;
	signal a0673 : integer;
	signal a0674 : integer;
	signal a0675 : integer;
	signal a0676 : integer;
	signal a0677 : integer;
	signal a0678 : integer;
	signal a0679 : integer;
	signal a0680 : integer;
	signal a0681 : integer;
	signal a0682 : integer;
	signal a0683 : integer;
	signal a0684 : integer;
	signal a0685 : integer;
	signal a0686 : integer;
	signal a0687 : integer;
	signal a0688 : integer;
	signal a0689 : integer;
	signal a0690 : integer;
	signal a0691 : integer;
	signal a0692 : integer;
	signal a0693 : integer;
	signal a0694 : integer;
	signal a0695 : integer;
	signal a0696 : integer;
	signal a0697 : integer;
	signal a0698 : integer;
	signal a0699 : integer;
	signal a0700 : integer;
	signal a0701 : integer;
	signal a0702 : integer;
	signal a0703 : integer;
	signal a0704 : integer;
	signal a0705 : integer;
	signal a0706 : integer;
	signal a0707 : integer;
	signal a0708 : integer;
	signal a0709 : integer;
	signal a0710 : integer;
	signal a0711 : integer;
	signal a0712 : integer;
	signal a0713 : integer;
	signal a0714 : integer;
	signal a0715 : integer;
	signal a0716 : integer;
	signal a0717 : integer;
	signal a0718 : integer;
	signal a0719 : integer;
	signal a0720 : integer;
	signal a0721 : integer;
	signal a0722 : integer;
	signal a0723 : integer;
	signal a0724 : integer;
	signal a0725 : integer;
	signal a0726 : integer;
	signal a0727 : integer;
	signal a0728 : integer;
	signal a0729 : integer;
	signal a0730 : integer;
	signal a0731 : integer;
	signal a0732 : integer;
	signal a0733 : integer;
	signal a0734 : integer;
	signal a0735 : integer;
	signal a0736 : integer;
	signal a0737 : integer;
	signal a0738 : integer;
	signal a0739 : integer;
	signal a0740 : integer;
	signal a0741 : integer;
	signal a0742 : integer;
	signal a0743 : integer;
	signal a0744 : integer;
	signal a0745 : integer;
	signal a0746 : integer;
	signal a0747 : integer;
	signal a0748 : integer;
	signal a0749 : integer;
	signal a0750 : integer;
	signal a0751 : integer;
	signal a0752 : integer;
	signal a0753 : integer;
	signal a0754 : integer;
	signal a0755 : integer;
	signal a0756 : integer;
	signal a0757 : integer;
	signal a0758 : integer;
	signal a0759 : integer;
	signal a0760 : integer;
	signal a0761 : integer;
	signal a0762 : integer;
	signal a0763 : integer;
	signal a0764 : integer;
	signal a0765 : integer;
	signal a0766 : integer;
	signal a0767 : integer;
	signal a0768 : integer;
	signal a0769 : integer;
	signal a0770 : integer;
	signal a0771 : integer;
	signal a0772 : integer;
	signal a0773 : integer;
	signal a0774 : integer;
	signal a0775 : integer;
	signal a0776 : integer;
	signal a0777 : integer;
	signal a0778 : integer;
	signal a0779 : integer;
	signal a0780 : integer;
	signal a0781 : integer;
	signal a0782 : integer;
	signal a0783 : integer;
	signal a0784 : integer;
	signal a0785 : integer;
	signal a0786 : integer;
	signal a0787 : integer;
	signal a0788 : integer;
	signal a0789 : integer;
	signal a0790 : integer;
	signal a0791 : integer;
	signal a0792 : integer;
	signal a0793 : integer;
	signal a0794 : integer;
	signal a0795 : integer;
	signal a0796 : integer;
	signal a0797 : integer;
	signal a0798 : integer;
	signal a0799 : integer;
	signal a0800 : integer;
	signal a0801 : integer;
	signal a0802 : integer;
	signal a0803 : integer;
	signal a0804 : integer;
	signal a0805 : integer;
	signal a0806 : integer;
	signal a0807 : integer;
	signal a0808 : integer;
	signal a0809 : integer;
	signal a0810 : integer;
	signal a0811 : integer;
	signal a0812 : integer;
	signal a0813 : integer;
	signal a0814 : integer;
	signal a0815 : integer;
	signal a0816 : integer;
	signal a0817 : integer;
	signal a0818 : integer;
	signal a0819 : integer;
	signal a0820 : integer;
	signal a0821 : integer;
	signal a0822 : integer;
	signal a0823 : integer;
	signal a0824 : integer;
	signal a0825 : integer;
	signal a0826 : integer;
	signal a0827 : integer;
	signal a0828 : integer;
	signal a0829 : integer;
	signal a0830 : integer;
	signal a0831 : integer;
	signal a0832 : integer;
	signal a0833 : integer;
	signal a0834 : integer;
	signal a0835 : integer;
	signal a0836 : integer;
	signal a0837 : integer;
	signal a0838 : integer;
	signal a0839 : integer;
	signal a0840 : integer;
	signal a0841 : integer;
	signal a0842 : integer;
	signal a0843 : integer;
	signal a0844 : integer;
	signal a0845 : integer;
	signal a0846 : integer;
	signal a0847 : integer;
	signal a0848 : integer;
	signal a0849 : integer;
	signal a0850 : integer;
	signal a0851 : integer;
	signal a0852 : integer;
	signal a0853 : integer;
	signal a0854 : integer;
	signal a0855 : integer;
	signal a0856 : integer;
	signal a0857 : integer;
	signal a0858 : integer;
	signal a0859 : integer;
	signal a0860 : integer;
	signal a0861 : integer;
	signal a0862 : integer;
	signal a0863 : integer;
	signal a0864 : integer;
	signal a0865 : integer;
	signal a0866 : integer;
	signal a0867 : integer;
	signal a0868 : integer;
	signal a0869 : integer;
	signal a0870 : integer;
	signal a0871 : integer;
	signal a0872 : integer;
	signal a0873 : integer;
	signal a0874 : integer;
	signal a0875 : integer;
	signal a0876 : integer;
	signal a0877 : integer;
	signal a0878 : integer;
	signal a0879 : integer;
	signal a0880 : integer;
	signal a0881 : integer;
	signal a0882 : integer;
	signal a0883 : integer;
	signal a0884 : integer;
	signal a0885 : integer;
	signal a0886 : integer;
	signal a0887 : integer;
	signal a0888 : integer;
	signal a0889 : integer;
	signal a0890 : integer;
	signal a0891 : integer;
	signal a0892 : integer;
	signal a0893 : integer;
	signal a0894 : integer;
	signal a0895 : integer;
	signal a0896 : integer;
	signal a0897 : integer;
	signal a0898 : integer;
	signal a0899 : integer;
	signal a0900 : integer;
	signal a0901 : integer;
	signal a0902 : integer;
	signal a0903 : integer;
	signal a0904 : integer;
	signal a0905 : integer;
	signal a0906 : integer;
	signal a0907 : integer;
	signal a0908 : integer;
	signal a0909 : integer;
	signal a0910 : integer;
	signal a0911 : integer;
	signal a0912 : integer;
	signal a0913 : integer;
	signal a0914 : integer;
	signal a0915 : integer;
	signal a0916 : integer;
	signal a0917 : integer;
	signal a0918 : integer;
	signal a0919 : integer;
	signal a0920 : integer;
	signal a0921 : integer;
	signal a0922 : integer;
	signal a0923 : integer;
	signal a0924 : integer;
	signal a0925 : integer;
	signal a0926 : integer;
	signal a0927 : integer;
	signal a0928 : integer;
	signal a0929 : integer;
	signal a0930 : integer;
	signal a0931 : integer;
	signal a0932 : integer;
	signal a0933 : integer;
	signal a0934 : integer;
	signal a0935 : integer;
	signal a0936 : integer;
	signal a0937 : integer;
	signal a0938 : integer;
	signal a0939 : integer;
	signal a0940 : integer;
	signal a0941 : integer;
	signal a0942 : integer;
	signal a0943 : integer;
	signal a0944 : integer;
	signal a0945 : integer;
	signal a0946 : integer;
	signal a0947 : integer;
	signal a0948 : integer;
	signal a0949 : integer;
	signal a0950 : integer;
	signal a0951 : integer;
	signal a0952 : integer;
	signal a0953 : integer;
	signal a0954 : integer;
	signal a0955 : integer;
	signal a0956 : integer;
	signal a0957 : integer;
	signal a0958 : integer;
	signal a0959 : integer;
	signal a0960 : integer;
	signal a0961 : integer;
	signal a0962 : integer;
	signal a0963 : integer;
	signal a0964 : integer;
	signal a0965 : integer;
	signal a0966 : integer;
	signal a0967 : integer;
	signal a0968 : integer;
	signal a0969 : integer;
	signal a0970 : integer;
	signal a0971 : integer;
	signal a0972 : integer;
	signal a0973 : integer;
	signal a0974 : integer;
	signal a0975 : integer;
	signal a0976 : integer;
	signal a0977 : integer;
	signal a0978 : integer;
	signal a0979 : integer;
	signal a0980 : integer;
	signal a0981 : integer;
	signal a0982 : integer;
	signal a0983 : integer;
	signal a0984 : integer;
	signal a0985 : integer;
	signal a0986 : integer;
	signal a0987 : integer;
	signal a0988 : integer;
	signal a0989 : integer;
	signal a0990 : integer;
	signal a0991 : integer;
	signal a0992 : integer;
	signal a0993 : integer;
	signal a0994 : integer;
	signal a0995 : integer;
	signal a0996 : integer;
	signal a0997 : integer;
	signal a0998 : integer;
	signal a0999 : integer;
	signal a1000 : integer;
	-- }}}
begin

	main: process(clk)
--{{{
	begin
		a0001 <= clk;
		a0002 <= clk;
		a0003 <= clk;
		a0004 <= clk;
		a0005 <= clk;
		a0006 <= clk;
		a0007 <= clk;
		a0008 <= clk;
		a0009 <= clk;
		a0010 <= clk;
		a0011 <= clk;
		a0012 <= clk;
		a0013 <= clk;
		a0014 <= clk;
		a0015 <= clk;
		a0016 <= clk;
		a0017 <= clk;
		a0018 <= clk;
		a0019 <= clk;
		a0020 <= clk;
		a0021 <= clk;
		a0022 <= clk;
		a0023 <= clk;
		a0024 <= clk;
		a0025 <= clk;
		a0026 <= clk;
		a0027 <= clk;
		a0028 <= clk;
		a0029 <= clk;
		a0030 <= clk;
		a0031 <= clk;
		a0032 <= clk;
		a0033 <= clk;
		a0034 <= clk;
		a0035 <= clk;
		a0036 <= clk;
		a0037 <= clk;
		a0038 <= clk;
		a0039 <= clk;
		a0040 <= clk;
		a0041 <= clk;
		a0042 <= clk;
		a0043 <= clk;
		a0044 <= clk;
		a0045 <= clk;
		a0046 <= clk;
		a0047 <= clk;
		a0048 <= clk;
		a0049 <= clk;
		a0050 <= clk;
		a0051 <= clk;
		a0052 <= clk;
		a0053 <= clk;
		a0054 <= clk;
		a0055 <= clk;
		a0056 <= clk;
		a0057 <= clk;
		a0058 <= clk;
		a0059 <= clk;
		a0060 <= clk;
		a0061 <= clk;
		a0062 <= clk;
		a0063 <= clk;
		a0064 <= clk;
		a0065 <= clk;
		a0066 <= clk;
		a0067 <= clk;
		a0068 <= clk;
		a0069 <= clk;
		a0070 <= clk;
		a0071 <= clk;
		a0072 <= clk;
		a0073 <= clk;
		a0074 <= clk;
		a0075 <= clk;
		a0076 <= clk;
		a0077 <= clk;
		a0078 <= clk;
		a0079 <= clk;
		a0080 <= clk;
		a0081 <= clk;
		a0082 <= clk;
		a0083 <= clk;
		a0084 <= clk;
		a0085 <= clk;
		a0086 <= clk;
		a0087 <= clk;
		a0088 <= clk;
		a0089 <= clk;
		a0090 <= clk;
		a0091 <= clk;
		a0092 <= clk;
		a0093 <= clk;
		a0094 <= clk;
		a0095 <= clk;
		a0096 <= clk;
		a0097 <= clk;
		a0098 <= clk;
		a0099 <= clk;
		a0100 <= clk;
		a0101 <= clk;
		a0102 <= clk;
		a0103 <= clk;
		a0104 <= clk;
		a0105 <= clk;
		a0106 <= clk;
		a0107 <= clk;
		a0108 <= clk;
		a0109 <= clk;
		a0110 <= clk;
		a0111 <= clk;
		a0112 <= clk;
		a0113 <= clk;
		a0114 <= clk;
		a0115 <= clk;
		a0116 <= clk;
		a0117 <= clk;
		a0118 <= clk;
		a0119 <= clk;
		a0120 <= clk;
		a0121 <= clk;
		a0122 <= clk;
		a0123 <= clk;
		a0124 <= clk;
		a0125 <= clk;
		a0126 <= clk;
		a0127 <= clk;
		a0128 <= clk;
		a0129 <= clk;
		a0130 <= clk;
		a0131 <= clk;
		a0132 <= clk;
		a0133 <= clk;
		a0134 <= clk;
		a0135 <= clk;
		a0136 <= clk;
		a0137 <= clk;
		a0138 <= clk;
		a0139 <= clk;
		a0140 <= clk;
		a0141 <= clk;
		a0142 <= clk;
		a0143 <= clk;
		a0144 <= clk;
		a0145 <= clk;
		a0146 <= clk;
		a0147 <= clk;
		a0148 <= clk;
		a0149 <= clk;
		a0150 <= clk;
		a0151 <= clk;
		a0152 <= clk;
		a0153 <= clk;
		a0154 <= clk;
		a0155 <= clk;
		a0156 <= clk;
		a0157 <= clk;
		a0158 <= clk;
		a0159 <= clk;
		a0160 <= clk;
		a0161 <= clk;
		a0162 <= clk;
		a0163 <= clk;
		a0164 <= clk;
		a0165 <= clk;
		a0166 <= clk;
		a0167 <= clk;
		a0168 <= clk;
		a0169 <= clk;
		a0170 <= clk;
		a0171 <= clk;
		a0172 <= clk;
		a0173 <= clk;
		a0174 <= clk;
		a0175 <= clk;
		a0176 <= clk;
		a0177 <= clk;
		a0178 <= clk;
		a0179 <= clk;
		a0180 <= clk;
		a0181 <= clk;
		a0182 <= clk;
		a0183 <= clk;
		a0184 <= clk;
		a0185 <= clk;
		a0186 <= clk;
		a0187 <= clk;
		a0188 <= clk;
		a0189 <= clk;
		a0190 <= clk;
		a0191 <= clk;
		a0192 <= clk;
		a0193 <= clk;
		a0194 <= clk;
		a0195 <= clk;
		a0196 <= clk;
		a0197 <= clk;
		a0198 <= clk;
		a0199 <= clk;
		a0200 <= clk;
		a0201 <= clk;
		a0202 <= clk;
		a0203 <= clk;
		a0204 <= clk;
		a0205 <= clk;
		a0206 <= clk;
		a0207 <= clk;
		a0208 <= clk;
		a0209 <= clk;
		a0210 <= clk;
		a0211 <= clk;
		a0212 <= clk;
		a0213 <= clk;
		a0214 <= clk;
		a0215 <= clk;
		a0216 <= clk;
		a0217 <= clk;
		a0218 <= clk;
		a0219 <= clk;
		a0220 <= clk;
		a0221 <= clk;
		a0222 <= clk;
		a0223 <= clk;
		a0224 <= clk;
		a0225 <= clk;
		a0226 <= clk;
		a0227 <= clk;
		a0228 <= clk;
		a0229 <= clk;
		a0230 <= clk;
		a0231 <= clk;
		a0232 <= clk;
		a0233 <= clk;
		a0234 <= clk;
		a0235 <= clk;
		a0236 <= clk;
		a0237 <= clk;
		a0238 <= clk;
		a0239 <= clk;
		a0240 <= clk;
		a0241 <= clk;
		a0242 <= clk;
		a0243 <= clk;
		a0244 <= clk;
		a0245 <= clk;
		a0246 <= clk;
		a0247 <= clk;
		a0248 <= clk;
		a0249 <= clk;
		a0250 <= clk;
		a0251 <= clk;
		a0252 <= clk;
		a0253 <= clk;
		a0254 <= clk;
		a0255 <= clk;
		a0256 <= clk;
		a0257 <= clk;
		a0258 <= clk;
		a0259 <= clk;
		a0260 <= clk;
		a0261 <= clk;
		a0262 <= clk;
		a0263 <= clk;
		a0264 <= clk;
		a0265 <= clk;
		a0266 <= clk;
		a0267 <= clk;
		a0268 <= clk;
		a0269 <= clk;
		a0270 <= clk;
		a0271 <= clk;
		a0272 <= clk;
		a0273 <= clk;
		a0274 <= clk;
		a0275 <= clk;
		a0276 <= clk;
		a0277 <= clk;
		a0278 <= clk;
		a0279 <= clk;
		a0280 <= clk;
		a0281 <= clk;
		a0282 <= clk;
		a0283 <= clk;
		a0284 <= clk;
		a0285 <= clk;
		a0286 <= clk;
		a0287 <= clk;
		a0288 <= clk;
		a0289 <= clk;
		a0290 <= clk;
		a0291 <= clk;
		a0292 <= clk;
		a0293 <= clk;
		a0294 <= clk;
		a0295 <= clk;
		a0296 <= clk;
		a0297 <= clk;
		a0298 <= clk;
		a0299 <= clk;
		a0300 <= clk;
		a0301 <= clk;
		a0302 <= clk;
		a0303 <= clk;
		a0304 <= clk;
		a0305 <= clk;
		a0306 <= clk;
		a0307 <= clk;
		a0308 <= clk;
		a0309 <= clk;
		a0310 <= clk;
		a0311 <= clk;
		a0312 <= clk;
		a0313 <= clk;
		a0314 <= clk;
		a0315 <= clk;
		a0316 <= clk;
		a0317 <= clk;
		a0318 <= clk;
		a0319 <= clk;
		a0320 <= clk;
		a0321 <= clk;
		a0322 <= clk;
		a0323 <= clk;
		a0324 <= clk;
		a0325 <= clk;
		a0326 <= clk;
		a0327 <= clk;
		a0328 <= clk;
		a0329 <= clk;
		a0330 <= clk;
		a0331 <= clk;
		a0332 <= clk;
		a0333 <= clk;
		a0334 <= clk;
		a0335 <= clk;
		a0336 <= clk;
		a0337 <= clk;
		a0338 <= clk;
		a0339 <= clk;
		a0340 <= clk;
		a0341 <= clk;
		a0342 <= clk;
		a0343 <= clk;
		a0344 <= clk;
		a0345 <= clk;
		a0346 <= clk;
		a0347 <= clk;
		a0348 <= clk;
		a0349 <= clk;
		a0350 <= clk;
		a0351 <= clk;
		a0352 <= clk;
		a0353 <= clk;
		a0354 <= clk;
		a0355 <= clk;
		a0356 <= clk;
		a0357 <= clk;
		a0358 <= clk;
		a0359 <= clk;
		a0360 <= clk;
		a0361 <= clk;
		a0362 <= clk;
		a0363 <= clk;
		a0364 <= clk;
		a0365 <= clk;
		a0366 <= clk;
		a0367 <= clk;
		a0368 <= clk;
		a0369 <= clk;
		a0370 <= clk;
		a0371 <= clk;
		a0372 <= clk;
		a0373 <= clk;
		a0374 <= clk;
		a0375 <= clk;
		a0376 <= clk;
		a0377 <= clk;
		a0378 <= clk;
		a0379 <= clk;
		a0380 <= clk;
		a0381 <= clk;
		a0382 <= clk;
		a0383 <= clk;
		a0384 <= clk;
		a0385 <= clk;
		a0386 <= clk;
		a0387 <= clk;
		a0388 <= clk;
		a0389 <= clk;
		a0390 <= clk;
		a0391 <= clk;
		a0392 <= clk;
		a0393 <= clk;
		a0394 <= clk;
		a0395 <= clk;
		a0396 <= clk;
		a0397 <= clk;
		a0398 <= clk;
		a0399 <= clk;
		a0400 <= clk;
		a0401 <= clk;
		a0402 <= clk;
		a0403 <= clk;
		a0404 <= clk;
		a0405 <= clk;
		a0406 <= clk;
		a0407 <= clk;
		a0408 <= clk;
		a0409 <= clk;
		a0410 <= clk;
		a0411 <= clk;
		a0412 <= clk;
		a0413 <= clk;
		a0414 <= clk;
		a0415 <= clk;
		a0416 <= clk;
		a0417 <= clk;
		a0418 <= clk;
		a0419 <= clk;
		a0420 <= clk;
		a0421 <= clk;
		a0422 <= clk;
		a0423 <= clk;
		a0424 <= clk;
		a0425 <= clk;
		a0426 <= clk;
		a0427 <= clk;
		a0428 <= clk;
		a0429 <= clk;
		a0430 <= clk;
		a0431 <= clk;
		a0432 <= clk;
		a0433 <= clk;
		a0434 <= clk;
		a0435 <= clk;
		a0436 <= clk;
		a0437 <= clk;
		a0438 <= clk;
		a0439 <= clk;
		a0440 <= clk;
		a0441 <= clk;
		a0442 <= clk;
		a0443 <= clk;
		a0444 <= clk;
		a0445 <= clk;
		a0446 <= clk;
		a0447 <= clk;
		a0448 <= clk;
		a0449 <= clk;
		a0450 <= clk;
		a0451 <= clk;
		a0452 <= clk;
		a0453 <= clk;
		a0454 <= clk;
		a0455 <= clk;
		a0456 <= clk;
		a0457 <= clk;
		a0458 <= clk;
		a0459 <= clk;
		a0460 <= clk;
		a0461 <= clk;
		a0462 <= clk;
		a0463 <= clk;
		a0464 <= clk;
		a0465 <= clk;
		a0466 <= clk;
		a0467 <= clk;
		a0468 <= clk;
		a0469 <= clk;
		a0470 <= clk;
		a0471 <= clk;
		a0472 <= clk;
		a0473 <= clk;
		a0474 <= clk;
		a0475 <= clk;
		a0476 <= clk;
		a0477 <= clk;
		a0478 <= clk;
		a0479 <= clk;
		a0480 <= clk;
		a0481 <= clk;
		a0482 <= clk;
		a0483 <= clk;
		a0484 <= clk;
		a0485 <= clk;
		a0486 <= clk;
		a0487 <= clk;
		a0488 <= clk;
		a0489 <= clk;
		a0490 <= clk;
		a0491 <= clk;
		a0492 <= clk;
		a0493 <= clk;
		a0494 <= clk;
		a0495 <= clk;
		a0496 <= clk;
		a0497 <= clk;
		a0498 <= clk;
		a0499 <= clk;
		a0500 <= clk;
		a0501 <= clk;
		a0502 <= clk;
		a0503 <= clk;
		a0504 <= clk;
		a0505 <= clk;
		a0506 <= clk;
		a0507 <= clk;
		a0508 <= clk;
		a0509 <= clk;
		a0510 <= clk;
		a0511 <= clk;
		a0512 <= clk;
		a0513 <= clk;
		a0514 <= clk;
		a0515 <= clk;
		a0516 <= clk;
		a0517 <= clk;
		a0518 <= clk;
		a0519 <= clk;
		a0520 <= clk;
		a0521 <= clk;
		a0522 <= clk;
		a0523 <= clk;
		a0524 <= clk;
		a0525 <= clk;
		a0526 <= clk;
		a0527 <= clk;
		a0528 <= clk;
		a0529 <= clk;
		a0530 <= clk;
		a0531 <= clk;
		a0532 <= clk;
		a0533 <= clk;
		a0534 <= clk;
		a0535 <= clk;
		a0536 <= clk;
		a0537 <= clk;
		a0538 <= clk;
		a0539 <= clk;
		a0540 <= clk;
		a0541 <= clk;
		a0542 <= clk;
		a0543 <= clk;
		a0544 <= clk;
		a0545 <= clk;
		a0546 <= clk;
		a0547 <= clk;
		a0548 <= clk;
		a0549 <= clk;
		a0550 <= clk;
		a0551 <= clk;
		a0552 <= clk;
		a0553 <= clk;
		a0554 <= clk;
		a0555 <= clk;
		a0556 <= clk;
		a0557 <= clk;
		a0558 <= clk;
		a0559 <= clk;
		a0560 <= clk;
		a0561 <= clk;
		a0562 <= clk;
		a0563 <= clk;
		a0564 <= clk;
		a0565 <= clk;
		a0566 <= clk;
		a0567 <= clk;
		a0568 <= clk;
		a0569 <= clk;
		a0570 <= clk;
		a0571 <= clk;
		a0572 <= clk;
		a0573 <= clk;
		a0574 <= clk;
		a0575 <= clk;
		a0576 <= clk;
		a0577 <= clk;
		a0578 <= clk;
		a0579 <= clk;
		a0580 <= clk;
		a0581 <= clk;
		a0582 <= clk;
		a0583 <= clk;
		a0584 <= clk;
		a0585 <= clk;
		a0586 <= clk;
		a0587 <= clk;
		a0588 <= clk;
		a0589 <= clk;
		a0590 <= clk;
		a0591 <= clk;
		a0592 <= clk;
		a0593 <= clk;
		a0594 <= clk;
		a0595 <= clk;
		a0596 <= clk;
		a0597 <= clk;
		a0598 <= clk;
		a0599 <= clk;
		a0600 <= clk;
		a0601 <= clk;
		a0602 <= clk;
		a0603 <= clk;
		a0604 <= clk;
		a0605 <= clk;
		a0606 <= clk;
		a0607 <= clk;
		a0608 <= clk;
		a0609 <= clk;
		a0610 <= clk;
		a0611 <= clk;
		a0612 <= clk;
		a0613 <= clk;
		a0614 <= clk;
		a0615 <= clk;
		a0616 <= clk;
		a0617 <= clk;
		a0618 <= clk;
		a0619 <= clk;
		a0620 <= clk;
		a0621 <= clk;
		a0622 <= clk;
		a0623 <= clk;
		a0624 <= clk;
		a0625 <= clk;
		a0626 <= clk;
		a0627 <= clk;
		a0628 <= clk;
		a0629 <= clk;
		a0630 <= clk;
		a0631 <= clk;
		a0632 <= clk;
		a0633 <= clk;
		a0634 <= clk;
		a0635 <= clk;
		a0636 <= clk;
		a0637 <= clk;
		a0638 <= clk;
		a0639 <= clk;
		a0640 <= clk;
		a0641 <= clk;
		a0642 <= clk;
		a0643 <= clk;
		a0644 <= clk;
		a0645 <= clk;
		a0646 <= clk;
		a0647 <= clk;
		a0648 <= clk;
		a0649 <= clk;
		a0650 <= clk;
		a0651 <= clk;
		a0652 <= clk;
		a0653 <= clk;
		a0654 <= clk;
		a0655 <= clk;
		a0656 <= clk;
		a0657 <= clk;
		a0658 <= clk;
		a0659 <= clk;
		a0660 <= clk;
		a0661 <= clk;
		a0662 <= clk;
		a0663 <= clk;
		a0664 <= clk;
		a0665 <= clk;
		a0666 <= clk;
		a0667 <= clk;
		a0668 <= clk;
		a0669 <= clk;
		a0670 <= clk;
		a0671 <= clk;
		a0672 <= clk;
		a0673 <= clk;
		a0674 <= clk;
		a0675 <= clk;
		a0676 <= clk;
		a0677 <= clk;
		a0678 <= clk;
		a0679 <= clk;
		a0680 <= clk;
		a0681 <= clk;
		a0682 <= clk;
		a0683 <= clk;
		a0684 <= clk;
		a0685 <= clk;
		a0686 <= clk;
		a0687 <= clk;
		a0688 <= clk;
		a0689 <= clk;
		a0690 <= clk;
		a0691 <= clk;
		a0692 <= clk;
		a0693 <= clk;
		a0694 <= clk;
		a0695 <= clk;
		a0696 <= clk;
		a0697 <= clk;
		a0698 <= clk;
		a0699 <= clk;
		a0700 <= clk;
		a0701 <= clk;
		a0702 <= clk;
		a0703 <= clk;
		a0704 <= clk;
		a0705 <= clk;
		a0706 <= clk;
		a0707 <= clk;
		a0708 <= clk;
		a0709 <= clk;
		a0710 <= clk;
		a0711 <= clk;
		a0712 <= clk;
		a0713 <= clk;
		a0714 <= clk;
		a0715 <= clk;
		a0716 <= clk;
		a0717 <= clk;
		a0718 <= clk;
		a0719 <= clk;
		a0720 <= clk;
		a0721 <= clk;
		a0722 <= clk;
		a0723 <= clk;
		a0724 <= clk;
		a0725 <= clk;
		a0726 <= clk;
		a0727 <= clk;
		a0728 <= clk;
		a0729 <= clk;
		a0730 <= clk;
		a0731 <= clk;
		a0732 <= clk;
		a0733 <= clk;
		a0734 <= clk;
		a0735 <= clk;
		a0736 <= clk;
		a0737 <= clk;
		a0738 <= clk;
		a0739 <= clk;
		a0740 <= clk;
		a0741 <= clk;
		a0742 <= clk;
		a0743 <= clk;
		a0744 <= clk;
		a0745 <= clk;
		a0746 <= clk;
		a0747 <= clk;
		a0748 <= clk;
		a0749 <= clk;
		a0750 <= clk;
		a0751 <= clk;
		a0752 <= clk;
		a0753 <= clk;
		a0754 <= clk;
		a0755 <= clk;
		a0756 <= clk;
		a0757 <= clk;
		a0758 <= clk;
		a0759 <= clk;
		a0760 <= clk;
		a0761 <= clk;
		a0762 <= clk;
		a0763 <= clk;
		a0764 <= clk;
		a0765 <= clk;
		a0766 <= clk;
		a0767 <= clk;
		a0768 <= clk;
		a0769 <= clk;
		a0770 <= clk;
		a0771 <= clk;
		a0772 <= clk;
		a0773 <= clk;
		a0774 <= clk;
		a0775 <= clk;
		a0776 <= clk;
		a0777 <= clk;
		a0778 <= clk;
		a0779 <= clk;
		a0780 <= clk;
		a0781 <= clk;
		a0782 <= clk;
		a0783 <= clk;
		a0784 <= clk;
		a0785 <= clk;
		a0786 <= clk;
		a0787 <= clk;
		a0788 <= clk;
		a0789 <= clk;
		a0790 <= clk;
		a0791 <= clk;
		a0792 <= clk;
		a0793 <= clk;
		a0794 <= clk;
		a0795 <= clk;
		a0796 <= clk;
		a0797 <= clk;
		a0798 <= clk;
		a0799 <= clk;
		a0800 <= clk;
		a0801 <= clk;
		a0802 <= clk;
		a0803 <= clk;
		a0804 <= clk;
		a0805 <= clk;
		a0806 <= clk;
		a0807 <= clk;
		a0808 <= clk;
		a0809 <= clk;
		a0810 <= clk;
		a0811 <= clk;
		a0812 <= clk;
		a0813 <= clk;
		a0814 <= clk;
		a0815 <= clk;
		a0816 <= clk;
		a0817 <= clk;
		a0818 <= clk;
		a0819 <= clk;
		a0820 <= clk;
		a0821 <= clk;
		a0822 <= clk;
		a0823 <= clk;
		a0824 <= clk;
		a0825 <= clk;
		a0826 <= clk;
		a0827 <= clk;
		a0828 <= clk;
		a0829 <= clk;
		a0830 <= clk;
		a0831 <= clk;
		a0832 <= clk;
		a0833 <= clk;
		a0834 <= clk;
		a0835 <= clk;
		a0836 <= clk;
		a0837 <= clk;
		a0838 <= clk;
		a0839 <= clk;
		a0840 <= clk;
		a0841 <= clk;
		a0842 <= clk;
		a0843 <= clk;
		a0844 <= clk;
		a0845 <= clk;
		a0846 <= clk;
		a0847 <= clk;
		a0848 <= clk;
		a0849 <= clk;
		a0850 <= clk;
		a0851 <= clk;
		a0852 <= clk;
		a0853 <= clk;
		a0854 <= clk;
		a0855 <= clk;
		a0856 <= clk;
		a0857 <= clk;
		a0858 <= clk;
		a0859 <= clk;
		a0860 <= clk;
		a0861 <= clk;
		a0862 <= clk;
		a0863 <= clk;
		a0864 <= clk;
		a0865 <= clk;
		a0866 <= clk;
		a0867 <= clk;
		a0868 <= clk;
		a0869 <= clk;
		a0870 <= clk;
		a0871 <= clk;
		a0872 <= clk;
		a0873 <= clk;
		a0874 <= clk;
		a0875 <= clk;
		a0876 <= clk;
		a0877 <= clk;
		a0878 <= clk;
		a0879 <= clk;
		a0880 <= clk;
		a0881 <= clk;
		a0882 <= clk;
		a0883 <= clk;
		a0884 <= clk;
		a0885 <= clk;
		a0886 <= clk;
		a0887 <= clk;
		a0888 <= clk;
		a0889 <= clk;
		a0890 <= clk;
		a0891 <= clk;
		a0892 <= clk;
		a0893 <= clk;
		a0894 <= clk;
		a0895 <= clk;
		a0896 <= clk;
		a0897 <= clk;
		a0898 <= clk;
		a0899 <= clk;
		a0900 <= clk;
		a0901 <= clk;
		a0902 <= clk;
		a0903 <= clk;
		a0904 <= clk;
		a0905 <= clk;
		a0906 <= clk;
		a0907 <= clk;
		a0908 <= clk;
		a0909 <= clk;
		a0910 <= clk;
		a0911 <= clk;
		a0912 <= clk;
		a0913 <= clk;
		a0914 <= clk;
		a0915 <= clk;
		a0916 <= clk;
		a0917 <= clk;
		a0918 <= clk;
		a0919 <= clk;
		a0920 <= clk;
		a0921 <= clk;
		a0922 <= clk;
		a0923 <= clk;
		a0924 <= clk;
		a0925 <= clk;
		a0926 <= clk;
		a0927 <= clk;
		a0928 <= clk;
		a0929 <= clk;
		a0930 <= clk;
		a0931 <= clk;
		a0932 <= clk;
		a0933 <= clk;
		a0934 <= clk;
		a0935 <= clk;
		a0936 <= clk;
		a0937 <= clk;
		a0938 <= clk;
		a0939 <= clk;
		a0940 <= clk;
		a0941 <= clk;
		a0942 <= clk;
		a0943 <= clk;
		a0944 <= clk;
		a0945 <= clk;
		a0946 <= clk;
		a0947 <= clk;
		a0948 <= clk;
		a0949 <= clk;
		a0950 <= clk;
		a0951 <= clk;
		a0952 <= clk;
		a0953 <= clk;
		a0954 <= clk;
		a0955 <= clk;
		a0956 <= clk;
		a0957 <= clk;
		a0958 <= clk;
		a0959 <= clk;
		a0960 <= clk;
		a0961 <= clk;
		a0962 <= clk;
		a0963 <= clk;
		a0964 <= clk;
		a0965 <= clk;
		a0966 <= clk;
		a0967 <= clk;
		a0968 <= clk;
		a0969 <= clk;
		a0970 <= clk;
		a0971 <= clk;
		a0972 <= clk;
		a0973 <= clk;
		a0974 <= clk;
		a0975 <= clk;
		a0976 <= clk;
		a0977 <= clk;
		a0978 <= clk;
		a0979 <= clk;
		a0980 <= clk;
		a0981 <= clk;
		a0982 <= clk;
		a0983 <= clk;
		a0984 <= clk;
		a0985 <= clk;
		a0986 <= clk;
		a0987 <= clk;
		a0988 <= clk;
		a0989 <= clk;
		a0990 <= clk;
		a0991 <= clk;
		a0992 <= clk;
		a0993 <= clk;
		a0994 <= clk;
		a0995 <= clk;
		a0996 <= clk;
		a0997 <= clk;
		a0998 <= clk;
		a0999 <= clk;
		a1000 <= clk;
        report "tick";
--}}}
    end process;

	terminator : process(clk)
	begin
		if clk >= CYCLES then
			assert false report "end of simulation" severity failure;
		-- else
		-- 	report "tick";
		end if;
	end process;

	clk <= (clk+1) after 1 us;
end;
