entity ENT00001_Test_Bench is
end entity ENT00001_Test_Bench;

architecture arch of ENT00001_Test_Bench is
	signal clk : integer := 0;
	constant CYCLES : integer := 1000;
begin

	main: process(clk)
--{{{
		variable a0001 : integer;
		variable a0002 : integer;
		variable a0003 : integer;
		variable a0004 : integer;
		variable a0005 : integer;
		variable a0006 : integer;
		variable a0007 : integer;
		variable a0008 : integer;
		variable a0009 : integer;
		variable a0010 : integer;
		variable a0011 : integer;
		variable a0012 : integer;
		variable a0013 : integer;
		variable a0014 : integer;
		variable a0015 : integer;
		variable a0016 : integer;
		variable a0017 : integer;
		variable a0018 : integer;
		variable a0019 : integer;
		variable a0020 : integer;
		variable a0021 : integer;
		variable a0022 : integer;
		variable a0023 : integer;
		variable a0024 : integer;
		variable a0025 : integer;
		variable a0026 : integer;
		variable a0027 : integer;
		variable a0028 : integer;
		variable a0029 : integer;
		variable a0030 : integer;
		variable a0031 : integer;
		variable a0032 : integer;
		variable a0033 : integer;
		variable a0034 : integer;
		variable a0035 : integer;
		variable a0036 : integer;
		variable a0037 : integer;
		variable a0038 : integer;
		variable a0039 : integer;
		variable a0040 : integer;
		variable a0041 : integer;
		variable a0042 : integer;
		variable a0043 : integer;
		variable a0044 : integer;
		variable a0045 : integer;
		variable a0046 : integer;
		variable a0047 : integer;
		variable a0048 : integer;
		variable a0049 : integer;
		variable a0050 : integer;
		variable a0051 : integer;
		variable a0052 : integer;
		variable a0053 : integer;
		variable a0054 : integer;
		variable a0055 : integer;
		variable a0056 : integer;
		variable a0057 : integer;
		variable a0058 : integer;
		variable a0059 : integer;
		variable a0060 : integer;
		variable a0061 : integer;
		variable a0062 : integer;
		variable a0063 : integer;
		variable a0064 : integer;
		variable a0065 : integer;
		variable a0066 : integer;
		variable a0067 : integer;
		variable a0068 : integer;
		variable a0069 : integer;
		variable a0070 : integer;
		variable a0071 : integer;
		variable a0072 : integer;
		variable a0073 : integer;
		variable a0074 : integer;
		variable a0075 : integer;
		variable a0076 : integer;
		variable a0077 : integer;
		variable a0078 : integer;
		variable a0079 : integer;
		variable a0080 : integer;
		variable a0081 : integer;
		variable a0082 : integer;
		variable a0083 : integer;
		variable a0084 : integer;
		variable a0085 : integer;
		variable a0086 : integer;
		variable a0087 : integer;
		variable a0088 : integer;
		variable a0089 : integer;
		variable a0090 : integer;
		variable a0091 : integer;
		variable a0092 : integer;
		variable a0093 : integer;
		variable a0094 : integer;
		variable a0095 : integer;
		variable a0096 : integer;
		variable a0097 : integer;
		variable a0098 : integer;
		variable a0099 : integer;
		variable a0100 : integer;
		variable a0101 : integer;
		variable a0102 : integer;
		variable a0103 : integer;
		variable a0104 : integer;
		variable a0105 : integer;
		variable a0106 : integer;
		variable a0107 : integer;
		variable a0108 : integer;
		variable a0109 : integer;
		variable a0110 : integer;
		variable a0111 : integer;
		variable a0112 : integer;
		variable a0113 : integer;
		variable a0114 : integer;
		variable a0115 : integer;
		variable a0116 : integer;
		variable a0117 : integer;
		variable a0118 : integer;
		variable a0119 : integer;
		variable a0120 : integer;
		variable a0121 : integer;
		variable a0122 : integer;
		variable a0123 : integer;
		variable a0124 : integer;
		variable a0125 : integer;
		variable a0126 : integer;
		variable a0127 : integer;
		variable a0128 : integer;
		variable a0129 : integer;
		variable a0130 : integer;
		variable a0131 : integer;
		variable a0132 : integer;
		variable a0133 : integer;
		variable a0134 : integer;
		variable a0135 : integer;
		variable a0136 : integer;
		variable a0137 : integer;
		variable a0138 : integer;
		variable a0139 : integer;
		variable a0140 : integer;
		variable a0141 : integer;
		variable a0142 : integer;
		variable a0143 : integer;
		variable a0144 : integer;
		variable a0145 : integer;
		variable a0146 : integer;
		variable a0147 : integer;
		variable a0148 : integer;
		variable a0149 : integer;
		variable a0150 : integer;
		variable a0151 : integer;
		variable a0152 : integer;
		variable a0153 : integer;
		variable a0154 : integer;
		variable a0155 : integer;
		variable a0156 : integer;
		variable a0157 : integer;
		variable a0158 : integer;
		variable a0159 : integer;
		variable a0160 : integer;
		variable a0161 : integer;
		variable a0162 : integer;
		variable a0163 : integer;
		variable a0164 : integer;
		variable a0165 : integer;
		variable a0166 : integer;
		variable a0167 : integer;
		variable a0168 : integer;
		variable a0169 : integer;
		variable a0170 : integer;
		variable a0171 : integer;
		variable a0172 : integer;
		variable a0173 : integer;
		variable a0174 : integer;
		variable a0175 : integer;
		variable a0176 : integer;
		variable a0177 : integer;
		variable a0178 : integer;
		variable a0179 : integer;
		variable a0180 : integer;
		variable a0181 : integer;
		variable a0182 : integer;
		variable a0183 : integer;
		variable a0184 : integer;
		variable a0185 : integer;
		variable a0186 : integer;
		variable a0187 : integer;
		variable a0188 : integer;
		variable a0189 : integer;
		variable a0190 : integer;
		variable a0191 : integer;
		variable a0192 : integer;
		variable a0193 : integer;
		variable a0194 : integer;
		variable a0195 : integer;
		variable a0196 : integer;
		variable a0197 : integer;
		variable a0198 : integer;
		variable a0199 : integer;
		variable a0200 : integer;
		variable a0201 : integer;
		variable a0202 : integer;
		variable a0203 : integer;
		variable a0204 : integer;
		variable a0205 : integer;
		variable a0206 : integer;
		variable a0207 : integer;
		variable a0208 : integer;
		variable a0209 : integer;
		variable a0210 : integer;
		variable a0211 : integer;
		variable a0212 : integer;
		variable a0213 : integer;
		variable a0214 : integer;
		variable a0215 : integer;
		variable a0216 : integer;
		variable a0217 : integer;
		variable a0218 : integer;
		variable a0219 : integer;
		variable a0220 : integer;
		variable a0221 : integer;
		variable a0222 : integer;
		variable a0223 : integer;
		variable a0224 : integer;
		variable a0225 : integer;
		variable a0226 : integer;
		variable a0227 : integer;
		variable a0228 : integer;
		variable a0229 : integer;
		variable a0230 : integer;
		variable a0231 : integer;
		variable a0232 : integer;
		variable a0233 : integer;
		variable a0234 : integer;
		variable a0235 : integer;
		variable a0236 : integer;
		variable a0237 : integer;
		variable a0238 : integer;
		variable a0239 : integer;
		variable a0240 : integer;
		variable a0241 : integer;
		variable a0242 : integer;
		variable a0243 : integer;
		variable a0244 : integer;
		variable a0245 : integer;
		variable a0246 : integer;
		variable a0247 : integer;
		variable a0248 : integer;
		variable a0249 : integer;
		variable a0250 : integer;
		variable a0251 : integer;
		variable a0252 : integer;
		variable a0253 : integer;
		variable a0254 : integer;
		variable a0255 : integer;
		variable a0256 : integer;
		variable a0257 : integer;
		variable a0258 : integer;
		variable a0259 : integer;
		variable a0260 : integer;
		variable a0261 : integer;
		variable a0262 : integer;
		variable a0263 : integer;
		variable a0264 : integer;
		variable a0265 : integer;
		variable a0266 : integer;
		variable a0267 : integer;
		variable a0268 : integer;
		variable a0269 : integer;
		variable a0270 : integer;
		variable a0271 : integer;
		variable a0272 : integer;
		variable a0273 : integer;
		variable a0274 : integer;
		variable a0275 : integer;
		variable a0276 : integer;
		variable a0277 : integer;
		variable a0278 : integer;
		variable a0279 : integer;
		variable a0280 : integer;
		variable a0281 : integer;
		variable a0282 : integer;
		variable a0283 : integer;
		variable a0284 : integer;
		variable a0285 : integer;
		variable a0286 : integer;
		variable a0287 : integer;
		variable a0288 : integer;
		variable a0289 : integer;
		variable a0290 : integer;
		variable a0291 : integer;
		variable a0292 : integer;
		variable a0293 : integer;
		variable a0294 : integer;
		variable a0295 : integer;
		variable a0296 : integer;
		variable a0297 : integer;
		variable a0298 : integer;
		variable a0299 : integer;
		variable a0300 : integer;
		variable a0301 : integer;
		variable a0302 : integer;
		variable a0303 : integer;
		variable a0304 : integer;
		variable a0305 : integer;
		variable a0306 : integer;
		variable a0307 : integer;
		variable a0308 : integer;
		variable a0309 : integer;
		variable a0310 : integer;
		variable a0311 : integer;
		variable a0312 : integer;
		variable a0313 : integer;
		variable a0314 : integer;
		variable a0315 : integer;
		variable a0316 : integer;
		variable a0317 : integer;
		variable a0318 : integer;
		variable a0319 : integer;
		variable a0320 : integer;
		variable a0321 : integer;
		variable a0322 : integer;
		variable a0323 : integer;
		variable a0324 : integer;
		variable a0325 : integer;
		variable a0326 : integer;
		variable a0327 : integer;
		variable a0328 : integer;
		variable a0329 : integer;
		variable a0330 : integer;
		variable a0331 : integer;
		variable a0332 : integer;
		variable a0333 : integer;
		variable a0334 : integer;
		variable a0335 : integer;
		variable a0336 : integer;
		variable a0337 : integer;
		variable a0338 : integer;
		variable a0339 : integer;
		variable a0340 : integer;
		variable a0341 : integer;
		variable a0342 : integer;
		variable a0343 : integer;
		variable a0344 : integer;
		variable a0345 : integer;
		variable a0346 : integer;
		variable a0347 : integer;
		variable a0348 : integer;
		variable a0349 : integer;
		variable a0350 : integer;
		variable a0351 : integer;
		variable a0352 : integer;
		variable a0353 : integer;
		variable a0354 : integer;
		variable a0355 : integer;
		variable a0356 : integer;
		variable a0357 : integer;
		variable a0358 : integer;
		variable a0359 : integer;
		variable a0360 : integer;
		variable a0361 : integer;
		variable a0362 : integer;
		variable a0363 : integer;
		variable a0364 : integer;
		variable a0365 : integer;
		variable a0366 : integer;
		variable a0367 : integer;
		variable a0368 : integer;
		variable a0369 : integer;
		variable a0370 : integer;
		variable a0371 : integer;
		variable a0372 : integer;
		variable a0373 : integer;
		variable a0374 : integer;
		variable a0375 : integer;
		variable a0376 : integer;
		variable a0377 : integer;
		variable a0378 : integer;
		variable a0379 : integer;
		variable a0380 : integer;
		variable a0381 : integer;
		variable a0382 : integer;
		variable a0383 : integer;
		variable a0384 : integer;
		variable a0385 : integer;
		variable a0386 : integer;
		variable a0387 : integer;
		variable a0388 : integer;
		variable a0389 : integer;
		variable a0390 : integer;
		variable a0391 : integer;
		variable a0392 : integer;
		variable a0393 : integer;
		variable a0394 : integer;
		variable a0395 : integer;
		variable a0396 : integer;
		variable a0397 : integer;
		variable a0398 : integer;
		variable a0399 : integer;
		variable a0400 : integer;
		variable a0401 : integer;
		variable a0402 : integer;
		variable a0403 : integer;
		variable a0404 : integer;
		variable a0405 : integer;
		variable a0406 : integer;
		variable a0407 : integer;
		variable a0408 : integer;
		variable a0409 : integer;
		variable a0410 : integer;
		variable a0411 : integer;
		variable a0412 : integer;
		variable a0413 : integer;
		variable a0414 : integer;
		variable a0415 : integer;
		variable a0416 : integer;
		variable a0417 : integer;
		variable a0418 : integer;
		variable a0419 : integer;
		variable a0420 : integer;
		variable a0421 : integer;
		variable a0422 : integer;
		variable a0423 : integer;
		variable a0424 : integer;
		variable a0425 : integer;
		variable a0426 : integer;
		variable a0427 : integer;
		variable a0428 : integer;
		variable a0429 : integer;
		variable a0430 : integer;
		variable a0431 : integer;
		variable a0432 : integer;
		variable a0433 : integer;
		variable a0434 : integer;
		variable a0435 : integer;
		variable a0436 : integer;
		variable a0437 : integer;
		variable a0438 : integer;
		variable a0439 : integer;
		variable a0440 : integer;
		variable a0441 : integer;
		variable a0442 : integer;
		variable a0443 : integer;
		variable a0444 : integer;
		variable a0445 : integer;
		variable a0446 : integer;
		variable a0447 : integer;
		variable a0448 : integer;
		variable a0449 : integer;
		variable a0450 : integer;
		variable a0451 : integer;
		variable a0452 : integer;
		variable a0453 : integer;
		variable a0454 : integer;
		variable a0455 : integer;
		variable a0456 : integer;
		variable a0457 : integer;
		variable a0458 : integer;
		variable a0459 : integer;
		variable a0460 : integer;
		variable a0461 : integer;
		variable a0462 : integer;
		variable a0463 : integer;
		variable a0464 : integer;
		variable a0465 : integer;
		variable a0466 : integer;
		variable a0467 : integer;
		variable a0468 : integer;
		variable a0469 : integer;
		variable a0470 : integer;
		variable a0471 : integer;
		variable a0472 : integer;
		variable a0473 : integer;
		variable a0474 : integer;
		variable a0475 : integer;
		variable a0476 : integer;
		variable a0477 : integer;
		variable a0478 : integer;
		variable a0479 : integer;
		variable a0480 : integer;
		variable a0481 : integer;
		variable a0482 : integer;
		variable a0483 : integer;
		variable a0484 : integer;
		variable a0485 : integer;
		variable a0486 : integer;
		variable a0487 : integer;
		variable a0488 : integer;
		variable a0489 : integer;
		variable a0490 : integer;
		variable a0491 : integer;
		variable a0492 : integer;
		variable a0493 : integer;
		variable a0494 : integer;
		variable a0495 : integer;
		variable a0496 : integer;
		variable a0497 : integer;
		variable a0498 : integer;
		variable a0499 : integer;
		variable a0500 : integer;
		variable a0501 : integer;
		variable a0502 : integer;
		variable a0503 : integer;
		variable a0504 : integer;
		variable a0505 : integer;
		variable a0506 : integer;
		variable a0507 : integer;
		variable a0508 : integer;
		variable a0509 : integer;
		variable a0510 : integer;
		variable a0511 : integer;
		variable a0512 : integer;
		variable a0513 : integer;
		variable a0514 : integer;
		variable a0515 : integer;
		variable a0516 : integer;
		variable a0517 : integer;
		variable a0518 : integer;
		variable a0519 : integer;
		variable a0520 : integer;
		variable a0521 : integer;
		variable a0522 : integer;
		variable a0523 : integer;
		variable a0524 : integer;
		variable a0525 : integer;
		variable a0526 : integer;
		variable a0527 : integer;
		variable a0528 : integer;
		variable a0529 : integer;
		variable a0530 : integer;
		variable a0531 : integer;
		variable a0532 : integer;
		variable a0533 : integer;
		variable a0534 : integer;
		variable a0535 : integer;
		variable a0536 : integer;
		variable a0537 : integer;
		variable a0538 : integer;
		variable a0539 : integer;
		variable a0540 : integer;
		variable a0541 : integer;
		variable a0542 : integer;
		variable a0543 : integer;
		variable a0544 : integer;
		variable a0545 : integer;
		variable a0546 : integer;
		variable a0547 : integer;
		variable a0548 : integer;
		variable a0549 : integer;
		variable a0550 : integer;
		variable a0551 : integer;
		variable a0552 : integer;
		variable a0553 : integer;
		variable a0554 : integer;
		variable a0555 : integer;
		variable a0556 : integer;
		variable a0557 : integer;
		variable a0558 : integer;
		variable a0559 : integer;
		variable a0560 : integer;
		variable a0561 : integer;
		variable a0562 : integer;
		variable a0563 : integer;
		variable a0564 : integer;
		variable a0565 : integer;
		variable a0566 : integer;
		variable a0567 : integer;
		variable a0568 : integer;
		variable a0569 : integer;
		variable a0570 : integer;
		variable a0571 : integer;
		variable a0572 : integer;
		variable a0573 : integer;
		variable a0574 : integer;
		variable a0575 : integer;
		variable a0576 : integer;
		variable a0577 : integer;
		variable a0578 : integer;
		variable a0579 : integer;
		variable a0580 : integer;
		variable a0581 : integer;
		variable a0582 : integer;
		variable a0583 : integer;
		variable a0584 : integer;
		variable a0585 : integer;
		variable a0586 : integer;
		variable a0587 : integer;
		variable a0588 : integer;
		variable a0589 : integer;
		variable a0590 : integer;
		variable a0591 : integer;
		variable a0592 : integer;
		variable a0593 : integer;
		variable a0594 : integer;
		variable a0595 : integer;
		variable a0596 : integer;
		variable a0597 : integer;
		variable a0598 : integer;
		variable a0599 : integer;
		variable a0600 : integer;
		variable a0601 : integer;
		variable a0602 : integer;
		variable a0603 : integer;
		variable a0604 : integer;
		variable a0605 : integer;
		variable a0606 : integer;
		variable a0607 : integer;
		variable a0608 : integer;
		variable a0609 : integer;
		variable a0610 : integer;
		variable a0611 : integer;
		variable a0612 : integer;
		variable a0613 : integer;
		variable a0614 : integer;
		variable a0615 : integer;
		variable a0616 : integer;
		variable a0617 : integer;
		variable a0618 : integer;
		variable a0619 : integer;
		variable a0620 : integer;
		variable a0621 : integer;
		variable a0622 : integer;
		variable a0623 : integer;
		variable a0624 : integer;
		variable a0625 : integer;
		variable a0626 : integer;
		variable a0627 : integer;
		variable a0628 : integer;
		variable a0629 : integer;
		variable a0630 : integer;
		variable a0631 : integer;
		variable a0632 : integer;
		variable a0633 : integer;
		variable a0634 : integer;
		variable a0635 : integer;
		variable a0636 : integer;
		variable a0637 : integer;
		variable a0638 : integer;
		variable a0639 : integer;
		variable a0640 : integer;
		variable a0641 : integer;
		variable a0642 : integer;
		variable a0643 : integer;
		variable a0644 : integer;
		variable a0645 : integer;
		variable a0646 : integer;
		variable a0647 : integer;
		variable a0648 : integer;
		variable a0649 : integer;
		variable a0650 : integer;
		variable a0651 : integer;
		variable a0652 : integer;
		variable a0653 : integer;
		variable a0654 : integer;
		variable a0655 : integer;
		variable a0656 : integer;
		variable a0657 : integer;
		variable a0658 : integer;
		variable a0659 : integer;
		variable a0660 : integer;
		variable a0661 : integer;
		variable a0662 : integer;
		variable a0663 : integer;
		variable a0664 : integer;
		variable a0665 : integer;
		variable a0666 : integer;
		variable a0667 : integer;
		variable a0668 : integer;
		variable a0669 : integer;
		variable a0670 : integer;
		variable a0671 : integer;
		variable a0672 : integer;
		variable a0673 : integer;
		variable a0674 : integer;
		variable a0675 : integer;
		variable a0676 : integer;
		variable a0677 : integer;
		variable a0678 : integer;
		variable a0679 : integer;
		variable a0680 : integer;
		variable a0681 : integer;
		variable a0682 : integer;
		variable a0683 : integer;
		variable a0684 : integer;
		variable a0685 : integer;
		variable a0686 : integer;
		variable a0687 : integer;
		variable a0688 : integer;
		variable a0689 : integer;
		variable a0690 : integer;
		variable a0691 : integer;
		variable a0692 : integer;
		variable a0693 : integer;
		variable a0694 : integer;
		variable a0695 : integer;
		variable a0696 : integer;
		variable a0697 : integer;
		variable a0698 : integer;
		variable a0699 : integer;
		variable a0700 : integer;
		variable a0701 : integer;
		variable a0702 : integer;
		variable a0703 : integer;
		variable a0704 : integer;
		variable a0705 : integer;
		variable a0706 : integer;
		variable a0707 : integer;
		variable a0708 : integer;
		variable a0709 : integer;
		variable a0710 : integer;
		variable a0711 : integer;
		variable a0712 : integer;
		variable a0713 : integer;
		variable a0714 : integer;
		variable a0715 : integer;
		variable a0716 : integer;
		variable a0717 : integer;
		variable a0718 : integer;
		variable a0719 : integer;
		variable a0720 : integer;
		variable a0721 : integer;
		variable a0722 : integer;
		variable a0723 : integer;
		variable a0724 : integer;
		variable a0725 : integer;
		variable a0726 : integer;
		variable a0727 : integer;
		variable a0728 : integer;
		variable a0729 : integer;
		variable a0730 : integer;
		variable a0731 : integer;
		variable a0732 : integer;
		variable a0733 : integer;
		variable a0734 : integer;
		variable a0735 : integer;
		variable a0736 : integer;
		variable a0737 : integer;
		variable a0738 : integer;
		variable a0739 : integer;
		variable a0740 : integer;
		variable a0741 : integer;
		variable a0742 : integer;
		variable a0743 : integer;
		variable a0744 : integer;
		variable a0745 : integer;
		variable a0746 : integer;
		variable a0747 : integer;
		variable a0748 : integer;
		variable a0749 : integer;
		variable a0750 : integer;
		variable a0751 : integer;
		variable a0752 : integer;
		variable a0753 : integer;
		variable a0754 : integer;
		variable a0755 : integer;
		variable a0756 : integer;
		variable a0757 : integer;
		variable a0758 : integer;
		variable a0759 : integer;
		variable a0760 : integer;
		variable a0761 : integer;
		variable a0762 : integer;
		variable a0763 : integer;
		variable a0764 : integer;
		variable a0765 : integer;
		variable a0766 : integer;
		variable a0767 : integer;
		variable a0768 : integer;
		variable a0769 : integer;
		variable a0770 : integer;
		variable a0771 : integer;
		variable a0772 : integer;
		variable a0773 : integer;
		variable a0774 : integer;
		variable a0775 : integer;
		variable a0776 : integer;
		variable a0777 : integer;
		variable a0778 : integer;
		variable a0779 : integer;
		variable a0780 : integer;
		variable a0781 : integer;
		variable a0782 : integer;
		variable a0783 : integer;
		variable a0784 : integer;
		variable a0785 : integer;
		variable a0786 : integer;
		variable a0787 : integer;
		variable a0788 : integer;
		variable a0789 : integer;
		variable a0790 : integer;
		variable a0791 : integer;
		variable a0792 : integer;
		variable a0793 : integer;
		variable a0794 : integer;
		variable a0795 : integer;
		variable a0796 : integer;
		variable a0797 : integer;
		variable a0798 : integer;
		variable a0799 : integer;
		variable a0800 : integer;
		variable a0801 : integer;
		variable a0802 : integer;
		variable a0803 : integer;
		variable a0804 : integer;
		variable a0805 : integer;
		variable a0806 : integer;
		variable a0807 : integer;
		variable a0808 : integer;
		variable a0809 : integer;
		variable a0810 : integer;
		variable a0811 : integer;
		variable a0812 : integer;
		variable a0813 : integer;
		variable a0814 : integer;
		variable a0815 : integer;
		variable a0816 : integer;
		variable a0817 : integer;
		variable a0818 : integer;
		variable a0819 : integer;
		variable a0820 : integer;
		variable a0821 : integer;
		variable a0822 : integer;
		variable a0823 : integer;
		variable a0824 : integer;
		variable a0825 : integer;
		variable a0826 : integer;
		variable a0827 : integer;
		variable a0828 : integer;
		variable a0829 : integer;
		variable a0830 : integer;
		variable a0831 : integer;
		variable a0832 : integer;
		variable a0833 : integer;
		variable a0834 : integer;
		variable a0835 : integer;
		variable a0836 : integer;
		variable a0837 : integer;
		variable a0838 : integer;
		variable a0839 : integer;
		variable a0840 : integer;
		variable a0841 : integer;
		variable a0842 : integer;
		variable a0843 : integer;
		variable a0844 : integer;
		variable a0845 : integer;
		variable a0846 : integer;
		variable a0847 : integer;
		variable a0848 : integer;
		variable a0849 : integer;
		variable a0850 : integer;
		variable a0851 : integer;
		variable a0852 : integer;
		variable a0853 : integer;
		variable a0854 : integer;
		variable a0855 : integer;
		variable a0856 : integer;
		variable a0857 : integer;
		variable a0858 : integer;
		variable a0859 : integer;
		variable a0860 : integer;
		variable a0861 : integer;
		variable a0862 : integer;
		variable a0863 : integer;
		variable a0864 : integer;
		variable a0865 : integer;
		variable a0866 : integer;
		variable a0867 : integer;
		variable a0868 : integer;
		variable a0869 : integer;
		variable a0870 : integer;
		variable a0871 : integer;
		variable a0872 : integer;
		variable a0873 : integer;
		variable a0874 : integer;
		variable a0875 : integer;
		variable a0876 : integer;
		variable a0877 : integer;
		variable a0878 : integer;
		variable a0879 : integer;
		variable a0880 : integer;
		variable a0881 : integer;
		variable a0882 : integer;
		variable a0883 : integer;
		variable a0884 : integer;
		variable a0885 : integer;
		variable a0886 : integer;
		variable a0887 : integer;
		variable a0888 : integer;
		variable a0889 : integer;
		variable a0890 : integer;
		variable a0891 : integer;
		variable a0892 : integer;
		variable a0893 : integer;
		variable a0894 : integer;
		variable a0895 : integer;
		variable a0896 : integer;
		variable a0897 : integer;
		variable a0898 : integer;
		variable a0899 : integer;
		variable a0900 : integer;
		variable a0901 : integer;
		variable a0902 : integer;
		variable a0903 : integer;
		variable a0904 : integer;
		variable a0905 : integer;
		variable a0906 : integer;
		variable a0907 : integer;
		variable a0908 : integer;
		variable a0909 : integer;
		variable a0910 : integer;
		variable a0911 : integer;
		variable a0912 : integer;
		variable a0913 : integer;
		variable a0914 : integer;
		variable a0915 : integer;
		variable a0916 : integer;
		variable a0917 : integer;
		variable a0918 : integer;
		variable a0919 : integer;
		variable a0920 : integer;
		variable a0921 : integer;
		variable a0922 : integer;
		variable a0923 : integer;
		variable a0924 : integer;
		variable a0925 : integer;
		variable a0926 : integer;
		variable a0927 : integer;
		variable a0928 : integer;
		variable a0929 : integer;
		variable a0930 : integer;
		variable a0931 : integer;
		variable a0932 : integer;
		variable a0933 : integer;
		variable a0934 : integer;
		variable a0935 : integer;
		variable a0936 : integer;
		variable a0937 : integer;
		variable a0938 : integer;
		variable a0939 : integer;
		variable a0940 : integer;
		variable a0941 : integer;
		variable a0942 : integer;
		variable a0943 : integer;
		variable a0944 : integer;
		variable a0945 : integer;
		variable a0946 : integer;
		variable a0947 : integer;
		variable a0948 : integer;
		variable a0949 : integer;
		variable a0950 : integer;
		variable a0951 : integer;
		variable a0952 : integer;
		variable a0953 : integer;
		variable a0954 : integer;
		variable a0955 : integer;
		variable a0956 : integer;
		variable a0957 : integer;
		variable a0958 : integer;
		variable a0959 : integer;
		variable a0960 : integer;
		variable a0961 : integer;
		variable a0962 : integer;
		variable a0963 : integer;
		variable a0964 : integer;
		variable a0965 : integer;
		variable a0966 : integer;
		variable a0967 : integer;
		variable a0968 : integer;
		variable a0969 : integer;
		variable a0970 : integer;
		variable a0971 : integer;
		variable a0972 : integer;
		variable a0973 : integer;
		variable a0974 : integer;
		variable a0975 : integer;
		variable a0976 : integer;
		variable a0977 : integer;
		variable a0978 : integer;
		variable a0979 : integer;
		variable a0980 : integer;
		variable a0981 : integer;
		variable a0982 : integer;
		variable a0983 : integer;
		variable a0984 : integer;
		variable a0985 : integer;
		variable a0986 : integer;
		variable a0987 : integer;
		variable a0988 : integer;
		variable a0989 : integer;
		variable a0990 : integer;
		variable a0991 : integer;
		variable a0992 : integer;
		variable a0993 : integer;
		variable a0994 : integer;
		variable a0995 : integer;
		variable a0996 : integer;
		variable a0997 : integer;
		variable a0998 : integer;
		variable a0999 : integer;
		variable a1000 : integer;
	begin

		a0001 := 1;
		a0002 := 2;
		a0003 := 3;
		a0004 := 4;
		a0005 := 5;
		a0006 := 6;
		a0007 := 7;
		a0008 := 8;
		a0009 := 9;
		a0010 := 10;
		a0011 := 11;
		a0012 := 12;
		a0013 := 13;
		a0014 := 14;
		a0015 := 15;
		a0016 := 16;
		a0017 := 17;
		a0018 := 18;
		a0019 := 19;
		a0020 := 20;
		a0021 := 21;
		a0022 := 22;
		a0023 := 23;
		a0024 := 24;
		a0025 := 25;
		a0026 := 26;
		a0027 := 27;
		a0028 := 28;
		a0029 := 29;
		a0030 := 30;
		a0031 := 31;
		a0032 := 32;
		a0033 := 33;
		a0034 := 34;
		a0035 := 35;
		a0036 := 36;
		a0037 := 37;
		a0038 := 38;
		a0039 := 39;
		a0040 := 40;
		a0041 := 41;
		a0042 := 42;
		a0043 := 43;
		a0044 := 44;
		a0045 := 45;
		a0046 := 46;
		a0047 := 47;
		a0048 := 48;
		a0049 := 49;
		a0050 := 50;
		a0051 := 51;
		a0052 := 52;
		a0053 := 53;
		a0054 := 54;
		a0055 := 55;
		a0056 := 56;
		a0057 := 57;
		a0058 := 58;
		a0059 := 59;
		a0060 := 60;
		a0061 := 61;
		a0062 := 62;
		a0063 := 63;
		a0064 := 64;
		a0065 := 65;
		a0066 := 66;
		a0067 := 67;
		a0068 := 68;
		a0069 := 69;
		a0070 := 70;
		a0071 := 71;
		a0072 := 72;
		a0073 := 73;
		a0074 := 74;
		a0075 := 75;
		a0076 := 76;
		a0077 := 77;
		a0078 := 78;
		a0079 := 79;
		a0080 := 80;
		a0081 := 81;
		a0082 := 82;
		a0083 := 83;
		a0084 := 84;
		a0085 := 85;
		a0086 := 86;
		a0087 := 87;
		a0088 := 88;
		a0089 := 89;
		a0090 := 90;
		a0091 := 91;
		a0092 := 92;
		a0093 := 93;
		a0094 := 94;
		a0095 := 95;
		a0096 := 96;
		a0097 := 97;
		a0098 := 98;
		a0099 := 99;
		a0100 := 100;
		a0101 := 101;
		a0102 := 102;
		a0103 := 103;
		a0104 := 104;
		a0105 := 105;
		a0106 := 106;
		a0107 := 107;
		a0108 := 108;
		a0109 := 109;
		a0110 := 110;
		a0111 := 111;
		a0112 := 112;
		a0113 := 113;
		a0114 := 114;
		a0115 := 115;
		a0116 := 116;
		a0117 := 117;
		a0118 := 118;
		a0119 := 119;
		a0120 := 120;
		a0121 := 121;
		a0122 := 122;
		a0123 := 123;
		a0124 := 124;
		a0125 := 125;
		a0126 := 126;
		a0127 := 127;
		a0128 := 128;
		a0129 := 129;
		a0130 := 130;
		a0131 := 131;
		a0132 := 132;
		a0133 := 133;
		a0134 := 134;
		a0135 := 135;
		a0136 := 136;
		a0137 := 137;
		a0138 := 138;
		a0139 := 139;
		a0140 := 140;
		a0141 := 141;
		a0142 := 142;
		a0143 := 143;
		a0144 := 144;
		a0145 := 145;
		a0146 := 146;
		a0147 := 147;
		a0148 := 148;
		a0149 := 149;
		a0150 := 150;
		a0151 := 151;
		a0152 := 152;
		a0153 := 153;
		a0154 := 154;
		a0155 := 155;
		a0156 := 156;
		a0157 := 157;
		a0158 := 158;
		a0159 := 159;
		a0160 := 160;
		a0161 := 161;
		a0162 := 162;
		a0163 := 163;
		a0164 := 164;
		a0165 := 165;
		a0166 := 166;
		a0167 := 167;
		a0168 := 168;
		a0169 := 169;
		a0170 := 170;
		a0171 := 171;
		a0172 := 172;
		a0173 := 173;
		a0174 := 174;
		a0175 := 175;
		a0176 := 176;
		a0177 := 177;
		a0178 := 178;
		a0179 := 179;
		a0180 := 180;
		a0181 := 181;
		a0182 := 182;
		a0183 := 183;
		a0184 := 184;
		a0185 := 185;
		a0186 := 186;
		a0187 := 187;
		a0188 := 188;
		a0189 := 189;
		a0190 := 190;
		a0191 := 191;
		a0192 := 192;
		a0193 := 193;
		a0194 := 194;
		a0195 := 195;
		a0196 := 196;
		a0197 := 197;
		a0198 := 198;
		a0199 := 199;
		a0200 := 200;
		a0201 := 201;
		a0202 := 202;
		a0203 := 203;
		a0204 := 204;
		a0205 := 205;
		a0206 := 206;
		a0207 := 207;
		a0208 := 208;
		a0209 := 209;
		a0210 := 210;
		a0211 := 211;
		a0212 := 212;
		a0213 := 213;
		a0214 := 214;
		a0215 := 215;
		a0216 := 216;
		a0217 := 217;
		a0218 := 218;
		a0219 := 219;
		a0220 := 220;
		a0221 := 221;
		a0222 := 222;
		a0223 := 223;
		a0224 := 224;
		a0225 := 225;
		a0226 := 226;
		a0227 := 227;
		a0228 := 228;
		a0229 := 229;
		a0230 := 230;
		a0231 := 231;
		a0232 := 232;
		a0233 := 233;
		a0234 := 234;
		a0235 := 235;
		a0236 := 236;
		a0237 := 237;
		a0238 := 238;
		a0239 := 239;
		a0240 := 240;
		a0241 := 241;
		a0242 := 242;
		a0243 := 243;
		a0244 := 244;
		a0245 := 245;
		a0246 := 246;
		a0247 := 247;
		a0248 := 248;
		a0249 := 249;
		a0250 := 250;
		a0251 := 251;
		a0252 := 252;
		a0253 := 253;
		a0254 := 254;
		a0255 := 255;
		a0256 := 256;
		a0257 := 257;
		a0258 := 258;
		a0259 := 259;
		a0260 := 260;
		a0261 := 261;
		a0262 := 262;
		a0263 := 263;
		a0264 := 264;
		a0265 := 265;
		a0266 := 266;
		a0267 := 267;
		a0268 := 268;
		a0269 := 269;
		a0270 := 270;
		a0271 := 271;
		a0272 := 272;
		a0273 := 273;
		a0274 := 274;
		a0275 := 275;
		a0276 := 276;
		a0277 := 277;
		a0278 := 278;
		a0279 := 279;
		a0280 := 280;
		a0281 := 281;
		a0282 := 282;
		a0283 := 283;
		a0284 := 284;
		a0285 := 285;
		a0286 := 286;
		a0287 := 287;
		a0288 := 288;
		a0289 := 289;
		a0290 := 290;
		a0291 := 291;
		a0292 := 292;
		a0293 := 293;
		a0294 := 294;
		a0295 := 295;
		a0296 := 296;
		a0297 := 297;
		a0298 := 298;
		a0299 := 299;
		a0300 := 300;
		a0301 := 301;
		a0302 := 302;
		a0303 := 303;
		a0304 := 304;
		a0305 := 305;
		a0306 := 306;
		a0307 := 307;
		a0308 := 308;
		a0309 := 309;
		a0310 := 310;
		a0311 := 311;
		a0312 := 312;
		a0313 := 313;
		a0314 := 314;
		a0315 := 315;
		a0316 := 316;
		a0317 := 317;
		a0318 := 318;
		a0319 := 319;
		a0320 := 320;
		a0321 := 321;
		a0322 := 322;
		a0323 := 323;
		a0324 := 324;
		a0325 := 325;
		a0326 := 326;
		a0327 := 327;
		a0328 := 328;
		a0329 := 329;
		a0330 := 330;
		a0331 := 331;
		a0332 := 332;
		a0333 := 333;
		a0334 := 334;
		a0335 := 335;
		a0336 := 336;
		a0337 := 337;
		a0338 := 338;
		a0339 := 339;
		a0340 := 340;
		a0341 := 341;
		a0342 := 342;
		a0343 := 343;
		a0344 := 344;
		a0345 := 345;
		a0346 := 346;
		a0347 := 347;
		a0348 := 348;
		a0349 := 349;
		a0350 := 350;
		a0351 := 351;
		a0352 := 352;
		a0353 := 353;
		a0354 := 354;
		a0355 := 355;
		a0356 := 356;
		a0357 := 357;
		a0358 := 358;
		a0359 := 359;
		a0360 := 360;
		a0361 := 361;
		a0362 := 362;
		a0363 := 363;
		a0364 := 364;
		a0365 := 365;
		a0366 := 366;
		a0367 := 367;
		a0368 := 368;
		a0369 := 369;
		a0370 := 370;
		a0371 := 371;
		a0372 := 372;
		a0373 := 373;
		a0374 := 374;
		a0375 := 375;
		a0376 := 376;
		a0377 := 377;
		a0378 := 378;
		a0379 := 379;
		a0380 := 380;
		a0381 := 381;
		a0382 := 382;
		a0383 := 383;
		a0384 := 384;
		a0385 := 385;
		a0386 := 386;
		a0387 := 387;
		a0388 := 388;
		a0389 := 389;
		a0390 := 390;
		a0391 := 391;
		a0392 := 392;
		a0393 := 393;
		a0394 := 394;
		a0395 := 395;
		a0396 := 396;
		a0397 := 397;
		a0398 := 398;
		a0399 := 399;
		a0400 := 400;
		a0401 := 401;
		a0402 := 402;
		a0403 := 403;
		a0404 := 404;
		a0405 := 405;
		a0406 := 406;
		a0407 := 407;
		a0408 := 408;
		a0409 := 409;
		a0410 := 410;
		a0411 := 411;
		a0412 := 412;
		a0413 := 413;
		a0414 := 414;
		a0415 := 415;
		a0416 := 416;
		a0417 := 417;
		a0418 := 418;
		a0419 := 419;
		a0420 := 420;
		a0421 := 421;
		a0422 := 422;
		a0423 := 423;
		a0424 := 424;
		a0425 := 425;
		a0426 := 426;
		a0427 := 427;
		a0428 := 428;
		a0429 := 429;
		a0430 := 430;
		a0431 := 431;
		a0432 := 432;
		a0433 := 433;
		a0434 := 434;
		a0435 := 435;
		a0436 := 436;
		a0437 := 437;
		a0438 := 438;
		a0439 := 439;
		a0440 := 440;
		a0441 := 441;
		a0442 := 442;
		a0443 := 443;
		a0444 := 444;
		a0445 := 445;
		a0446 := 446;
		a0447 := 447;
		a0448 := 448;
		a0449 := 449;
		a0450 := 450;
		a0451 := 451;
		a0452 := 452;
		a0453 := 453;
		a0454 := 454;
		a0455 := 455;
		a0456 := 456;
		a0457 := 457;
		a0458 := 458;
		a0459 := 459;
		a0460 := 460;
		a0461 := 461;
		a0462 := 462;
		a0463 := 463;
		a0464 := 464;
		a0465 := 465;
		a0466 := 466;
		a0467 := 467;
		a0468 := 468;
		a0469 := 469;
		a0470 := 470;
		a0471 := 471;
		a0472 := 472;
		a0473 := 473;
		a0474 := 474;
		a0475 := 475;
		a0476 := 476;
		a0477 := 477;
		a0478 := 478;
		a0479 := 479;
		a0480 := 480;
		a0481 := 481;
		a0482 := 482;
		a0483 := 483;
		a0484 := 484;
		a0485 := 485;
		a0486 := 486;
		a0487 := 487;
		a0488 := 488;
		a0489 := 489;
		a0490 := 490;
		a0491 := 491;
		a0492 := 492;
		a0493 := 493;
		a0494 := 494;
		a0495 := 495;
		a0496 := 496;
		a0497 := 497;
		a0498 := 498;
		a0499 := 499;
		a0500 := 500;
		a0501 := 501;
		a0502 := 502;
		a0503 := 503;
		a0504 := 504;
		a0505 := 505;
		a0506 := 506;
		a0507 := 507;
		a0508 := 508;
		a0509 := 509;
		a0510 := 510;
		a0511 := 511;
		a0512 := 512;
		a0513 := 513;
		a0514 := 514;
		a0515 := 515;
		a0516 := 516;
		a0517 := 517;
		a0518 := 518;
		a0519 := 519;
		a0520 := 520;
		a0521 := 521;
		a0522 := 522;
		a0523 := 523;
		a0524 := 524;
		a0525 := 525;
		a0526 := 526;
		a0527 := 527;
		a0528 := 528;
		a0529 := 529;
		a0530 := 530;
		a0531 := 531;
		a0532 := 532;
		a0533 := 533;
		a0534 := 534;
		a0535 := 535;
		a0536 := 536;
		a0537 := 537;
		a0538 := 538;
		a0539 := 539;
		a0540 := 540;
		a0541 := 541;
		a0542 := 542;
		a0543 := 543;
		a0544 := 544;
		a0545 := 545;
		a0546 := 546;
		a0547 := 547;
		a0548 := 548;
		a0549 := 549;
		a0550 := 550;
		a0551 := 551;
		a0552 := 552;
		a0553 := 553;
		a0554 := 554;
		a0555 := 555;
		a0556 := 556;
		a0557 := 557;
		a0558 := 558;
		a0559 := 559;
		a0560 := 560;
		a0561 := 561;
		a0562 := 562;
		a0563 := 563;
		a0564 := 564;
		a0565 := 565;
		a0566 := 566;
		a0567 := 567;
		a0568 := 568;
		a0569 := 569;
		a0570 := 570;
		a0571 := 571;
		a0572 := 572;
		a0573 := 573;
		a0574 := 574;
		a0575 := 575;
		a0576 := 576;
		a0577 := 577;
		a0578 := 578;
		a0579 := 579;
		a0580 := 580;
		a0581 := 581;
		a0582 := 582;
		a0583 := 583;
		a0584 := 584;
		a0585 := 585;
		a0586 := 586;
		a0587 := 587;
		a0588 := 588;
		a0589 := 589;
		a0590 := 590;
		a0591 := 591;
		a0592 := 592;
		a0593 := 593;
		a0594 := 594;
		a0595 := 595;
		a0596 := 596;
		a0597 := 597;
		a0598 := 598;
		a0599 := 599;
		a0600 := 600;
		a0601 := 601;
		a0602 := 602;
		a0603 := 603;
		a0604 := 604;
		a0605 := 605;
		a0606 := 606;
		a0607 := 607;
		a0608 := 608;
		a0609 := 609;
		a0610 := 610;
		a0611 := 611;
		a0612 := 612;
		a0613 := 613;
		a0614 := 614;
		a0615 := 615;
		a0616 := 616;
		a0617 := 617;
		a0618 := 618;
		a0619 := 619;
		a0620 := 620;
		a0621 := 621;
		a0622 := 622;
		a0623 := 623;
		a0624 := 624;
		a0625 := 625;
		a0626 := 626;
		a0627 := 627;
		a0628 := 628;
		a0629 := 629;
		a0630 := 630;
		a0631 := 631;
		a0632 := 632;
		a0633 := 633;
		a0634 := 634;
		a0635 := 635;
		a0636 := 636;
		a0637 := 637;
		a0638 := 638;
		a0639 := 639;
		a0640 := 640;
		a0641 := 641;
		a0642 := 642;
		a0643 := 643;
		a0644 := 644;
		a0645 := 645;
		a0646 := 646;
		a0647 := 647;
		a0648 := 648;
		a0649 := 649;
		a0650 := 650;
		a0651 := 651;
		a0652 := 652;
		a0653 := 653;
		a0654 := 654;
		a0655 := 655;
		a0656 := 656;
		a0657 := 657;
		a0658 := 658;
		a0659 := 659;
		a0660 := 660;
		a0661 := 661;
		a0662 := 662;
		a0663 := 663;
		a0664 := 664;
		a0665 := 665;
		a0666 := 666;
		a0667 := 667;
		a0668 := 668;
		a0669 := 669;
		a0670 := 670;
		a0671 := 671;
		a0672 := 672;
		a0673 := 673;
		a0674 := 674;
		a0675 := 675;
		a0676 := 676;
		a0677 := 677;
		a0678 := 678;
		a0679 := 679;
		a0680 := 680;
		a0681 := 681;
		a0682 := 682;
		a0683 := 683;
		a0684 := 684;
		a0685 := 685;
		a0686 := 686;
		a0687 := 687;
		a0688 := 688;
		a0689 := 689;
		a0690 := 690;
		a0691 := 691;
		a0692 := 692;
		a0693 := 693;
		a0694 := 694;
		a0695 := 695;
		a0696 := 696;
		a0697 := 697;
		a0698 := 698;
		a0699 := 699;
		a0700 := 700;
		a0701 := 701;
		a0702 := 702;
		a0703 := 703;
		a0704 := 704;
		a0705 := 705;
		a0706 := 706;
		a0707 := 707;
		a0708 := 708;
		a0709 := 709;
		a0710 := 710;
		a0711 := 711;
		a0712 := 712;
		a0713 := 713;
		a0714 := 714;
		a0715 := 715;
		a0716 := 716;
		a0717 := 717;
		a0718 := 718;
		a0719 := 719;
		a0720 := 720;
		a0721 := 721;
		a0722 := 722;
		a0723 := 723;
		a0724 := 724;
		a0725 := 725;
		a0726 := 726;
		a0727 := 727;
		a0728 := 728;
		a0729 := 729;
		a0730 := 730;
		a0731 := 731;
		a0732 := 732;
		a0733 := 733;
		a0734 := 734;
		a0735 := 735;
		a0736 := 736;
		a0737 := 737;
		a0738 := 738;
		a0739 := 739;
		a0740 := 740;
		a0741 := 741;
		a0742 := 742;
		a0743 := 743;
		a0744 := 744;
		a0745 := 745;
		a0746 := 746;
		a0747 := 747;
		a0748 := 748;
		a0749 := 749;
		a0750 := 750;
		a0751 := 751;
		a0752 := 752;
		a0753 := 753;
		a0754 := 754;
		a0755 := 755;
		a0756 := 756;
		a0757 := 757;
		a0758 := 758;
		a0759 := 759;
		a0760 := 760;
		a0761 := 761;
		a0762 := 762;
		a0763 := 763;
		a0764 := 764;
		a0765 := 765;
		a0766 := 766;
		a0767 := 767;
		a0768 := 768;
		a0769 := 769;
		a0770 := 770;
		a0771 := 771;
		a0772 := 772;
		a0773 := 773;
		a0774 := 774;
		a0775 := 775;
		a0776 := 776;
		a0777 := 777;
		a0778 := 778;
		a0779 := 779;
		a0780 := 780;
		a0781 := 781;
		a0782 := 782;
		a0783 := 783;
		a0784 := 784;
		a0785 := 785;
		a0786 := 786;
		a0787 := 787;
		a0788 := 788;
		a0789 := 789;
		a0790 := 790;
		a0791 := 791;
		a0792 := 792;
		a0793 := 793;
		a0794 := 794;
		a0795 := 795;
		a0796 := 796;
		a0797 := 797;
		a0798 := 798;
		a0799 := 799;
		a0800 := 800;
		a0801 := 801;
		a0802 := 802;
		a0803 := 803;
		a0804 := 804;
		a0805 := 805;
		a0806 := 806;
		a0807 := 807;
		a0808 := 808;
		a0809 := 809;
		a0810 := 810;
		a0811 := 811;
		a0812 := 812;
		a0813 := 813;
		a0814 := 814;
		a0815 := 815;
		a0816 := 816;
		a0817 := 817;
		a0818 := 818;
		a0819 := 819;
		a0820 := 820;
		a0821 := 821;
		a0822 := 822;
		a0823 := 823;
		a0824 := 824;
		a0825 := 825;
		a0826 := 826;
		a0827 := 827;
		a0828 := 828;
		a0829 := 829;
		a0830 := 830;
		a0831 := 831;
		a0832 := 832;
		a0833 := 833;
		a0834 := 834;
		a0835 := 835;
		a0836 := 836;
		a0837 := 837;
		a0838 := 838;
		a0839 := 839;
		a0840 := 840;
		a0841 := 841;
		a0842 := 842;
		a0843 := 843;
		a0844 := 844;
		a0845 := 845;
		a0846 := 846;
		a0847 := 847;
		a0848 := 848;
		a0849 := 849;
		a0850 := 850;
		a0851 := 851;
		a0852 := 852;
		a0853 := 853;
		a0854 := 854;
		a0855 := 855;
		a0856 := 856;
		a0857 := 857;
		a0858 := 858;
		a0859 := 859;
		a0860 := 860;
		a0861 := 861;
		a0862 := 862;
		a0863 := 863;
		a0864 := 864;
		a0865 := 865;
		a0866 := 866;
		a0867 := 867;
		a0868 := 868;
		a0869 := 869;
		a0870 := 870;
		a0871 := 871;
		a0872 := 872;
		a0873 := 873;
		a0874 := 874;
		a0875 := 875;
		a0876 := 876;
		a0877 := 877;
		a0878 := 878;
		a0879 := 879;
		a0880 := 880;
		a0881 := 881;
		a0882 := 882;
		a0883 := 883;
		a0884 := 884;
		a0885 := 885;
		a0886 := 886;
		a0887 := 887;
		a0888 := 888;
		a0889 := 889;
		a0890 := 890;
		a0891 := 891;
		a0892 := 892;
		a0893 := 893;
		a0894 := 894;
		a0895 := 895;
		a0896 := 896;
		a0897 := 897;
		a0898 := 898;
		a0899 := 899;
		a0900 := 900;
		a0901 := 901;
		a0902 := 902;
		a0903 := 903;
		a0904 := 904;
		a0905 := 905;
		a0906 := 906;
		a0907 := 907;
		a0908 := 908;
		a0909 := 909;
		a0910 := 910;
		a0911 := 911;
		a0912 := 912;
		a0913 := 913;
		a0914 := 914;
		a0915 := 915;
		a0916 := 916;
		a0917 := 917;
		a0918 := 918;
		a0919 := 919;
		a0920 := 920;
		a0921 := 921;
		a0922 := 922;
		a0923 := 923;
		a0924 := 924;
		a0925 := 925;
		a0926 := 926;
		a0927 := 927;
		a0928 := 928;
		a0929 := 929;
		a0930 := 930;
		a0931 := 931;
		a0932 := 932;
		a0933 := 933;
		a0934 := 934;
		a0935 := 935;
		a0936 := 936;
		a0937 := 937;
		a0938 := 938;
		a0939 := 939;
		a0940 := 940;
		a0941 := 941;
		a0942 := 942;
		a0943 := 943;
		a0944 := 944;
		a0945 := 945;
		a0946 := 946;
		a0947 := 947;
		a0948 := 948;
		a0949 := 949;
		a0950 := 950;
		a0951 := 951;
		a0952 := 952;
		a0953 := 953;
		a0954 := 954;
		a0955 := 955;
		a0956 := 956;
		a0957 := 957;
		a0958 := 958;
		a0959 := 959;
		a0960 := 960;
		a0961 := 961;
		a0962 := 962;
		a0963 := 963;
		a0964 := 964;
		a0965 := 965;
		a0966 := 966;
		a0967 := 967;
		a0968 := 968;
		a0969 := 969;
		a0970 := 970;
		a0971 := 971;
		a0972 := 972;
		a0973 := 973;
		a0974 := 974;
		a0975 := 975;
		a0976 := 976;
		a0977 := 977;
		a0978 := 978;
		a0979 := 979;
		a0980 := 980;
		a0981 := 981;
		a0982 := 982;
		a0983 := 983;
		a0984 := 984;
		a0985 := 985;
		a0986 := 986;
		a0987 := 987;
		a0988 := 988;
		a0989 := 989;
		a0990 := 990;
		a0991 := 991;
		a0992 := 992;
		a0993 := 993;
		a0994 := 994;
		a0995 := 995;
		a0996 := 996;
		a0997 := 997;
		a0998 := 998;
		a0999 := 999;
		a1000 := 1000;
        -- report "tick";
--}}}
    end process;

	terminator : process(clk)
	begin
		if clk >= CYCLES then
			assert false report "end of simulation" severity failure;
		-- else
		-- 	report "tick";
		end if;
	end process;

	clk <= (clk+1) after 1 us;
end;
