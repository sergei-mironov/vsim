-- 500 variable assignments in 2 processes. Assigning a signal.

entity main is
end entity main ;

architecture arch of main is
	signal clk : integer := 0;
	constant CYCLES : integer := 1000;
begin

	main: process(clk)
		--{{{
		variable a0502 : integer;
		variable a0503 : integer;
		variable a0504 : integer;
		variable a0505 : integer;
		variable a0506 : integer;
		variable a0507 : integer;
		variable a0508 : integer;
		variable a0509 : integer;
		variable a0510 : integer;
		variable a0511 : integer;
		variable a0512 : integer;
		variable a0513 : integer;
		variable a0514 : integer;
		variable a0515 : integer;
		variable a0516 : integer;
		variable a0517 : integer;
		variable a0518 : integer;
		variable a0519 : integer;
		variable a0520 : integer;
		variable a0521 : integer;
		variable a0522 : integer;
		variable a0523 : integer;
		variable a0524 : integer;
		variable a0525 : integer;
		variable a0526 : integer;
		variable a0527 : integer;
		variable a0528 : integer;
		variable a0529 : integer;
		variable a0530 : integer;
		variable a0531 : integer;
		variable a0532 : integer;
		variable a0533 : integer;
		variable a0534 : integer;
		variable a0535 : integer;
		variable a0536 : integer;
		variable a0537 : integer;
		variable a0538 : integer;
		variable a0539 : integer;
		variable a0540 : integer;
		variable a0541 : integer;
		variable a0542 : integer;
		variable a0543 : integer;
		variable a0544 : integer;
		variable a0545 : integer;
		variable a0546 : integer;
		variable a0547 : integer;
		variable a0548 : integer;
		variable a0549 : integer;
		variable a0550 : integer;
		variable a0551 : integer;
		variable a0552 : integer;
		variable a0553 : integer;
		variable a0554 : integer;
		variable a0555 : integer;
		variable a0556 : integer;
		variable a0557 : integer;
		variable a0558 : integer;
		variable a0559 : integer;
		variable a0560 : integer;
		variable a0561 : integer;
		variable a0562 : integer;
		variable a0563 : integer;
		variable a0564 : integer;
		variable a0565 : integer;
		variable a0566 : integer;
		variable a0567 : integer;
		variable a0568 : integer;
		variable a0569 : integer;
		variable a0570 : integer;
		variable a0571 : integer;
		variable a0572 : integer;
		variable a0573 : integer;
		variable a0574 : integer;
		variable a0575 : integer;
		variable a0576 : integer;
		variable a0577 : integer;
		variable a0578 : integer;
		variable a0579 : integer;
		variable a0580 : integer;
		variable a0581 : integer;
		variable a0582 : integer;
		variable a0583 : integer;
		variable a0584 : integer;
		variable a0585 : integer;
		variable a0586 : integer;
		variable a0587 : integer;
		variable a0588 : integer;
		variable a0589 : integer;
		variable a0590 : integer;
		variable a0591 : integer;
		variable a0592 : integer;
		variable a0593 : integer;
		variable a0594 : integer;
		variable a0595 : integer;
		variable a0596 : integer;
		variable a0597 : integer;
		variable a0598 : integer;
		variable a0599 : integer;
		variable a0600 : integer;
		variable a0601 : integer;
		variable a0602 : integer;
		variable a0603 : integer;
		variable a0604 : integer;
		variable a0605 : integer;
		variable a0606 : integer;
		variable a0607 : integer;
		variable a0608 : integer;
		variable a0609 : integer;
		variable a0610 : integer;
		variable a0611 : integer;
		variable a0612 : integer;
		variable a0613 : integer;
		variable a0614 : integer;
		variable a0615 : integer;
		variable a0616 : integer;
		variable a0617 : integer;
		variable a0618 : integer;
		variable a0619 : integer;
		variable a0620 : integer;
		variable a0621 : integer;
		variable a0622 : integer;
		variable a0623 : integer;
		variable a0624 : integer;
		variable a0625 : integer;
		variable a0626 : integer;
		variable a0627 : integer;
		variable a0628 : integer;
		variable a0629 : integer;
		variable a0630 : integer;
		variable a0631 : integer;
		variable a0632 : integer;
		variable a0633 : integer;
		variable a0634 : integer;
		variable a0635 : integer;
		variable a0636 : integer;
		variable a0637 : integer;
		variable a0638 : integer;
		variable a0639 : integer;
		variable a0640 : integer;
		variable a0641 : integer;
		variable a0642 : integer;
		variable a0643 : integer;
		variable a0644 : integer;
		variable a0645 : integer;
		variable a0646 : integer;
		variable a0647 : integer;
		variable a0648 : integer;
		variable a0649 : integer;
		variable a0650 : integer;
		variable a0651 : integer;
		variable a0652 : integer;
		variable a0653 : integer;
		variable a0654 : integer;
		variable a0655 : integer;
		variable a0656 : integer;
		variable a0657 : integer;
		variable a0658 : integer;
		variable a0659 : integer;
		variable a0660 : integer;
		variable a0661 : integer;
		variable a0662 : integer;
		variable a0663 : integer;
		variable a0664 : integer;
		variable a0665 : integer;
		variable a0666 : integer;
		variable a0667 : integer;
		variable a0668 : integer;
		variable a0669 : integer;
		variable a0670 : integer;
		variable a0671 : integer;
		variable a0672 : integer;
		variable a0673 : integer;
		variable a0674 : integer;
		variable a0675 : integer;
		variable a0676 : integer;
		variable a0677 : integer;
		variable a0678 : integer;
		variable a0679 : integer;
		variable a0680 : integer;
		variable a0681 : integer;
		variable a0682 : integer;
		variable a0683 : integer;
		variable a0684 : integer;
		variable a0685 : integer;
		variable a0686 : integer;
		variable a0687 : integer;
		variable a0688 : integer;
		variable a0689 : integer;
		variable a0690 : integer;
		variable a0691 : integer;
		variable a0692 : integer;
		variable a0693 : integer;
		variable a0694 : integer;
		variable a0695 : integer;
		variable a0696 : integer;
		variable a0697 : integer;
		variable a0698 : integer;
		variable a0699 : integer;
		variable a0700 : integer;
		variable a0701 : integer;
		variable a0702 : integer;
		variable a0703 : integer;
		variable a0704 : integer;
		variable a0705 : integer;
		variable a0706 : integer;
		variable a0707 : integer;
		variable a0708 : integer;
		variable a0709 : integer;
		variable a0710 : integer;
		variable a0711 : integer;
		variable a0712 : integer;
		variable a0713 : integer;
		variable a0714 : integer;
		variable a0715 : integer;
		variable a0716 : integer;
		variable a0717 : integer;
		variable a0718 : integer;
		variable a0719 : integer;
		variable a0720 : integer;
		variable a0721 : integer;
		variable a0722 : integer;
		variable a0723 : integer;
		variable a0724 : integer;
		variable a0725 : integer;
		variable a0726 : integer;
		variable a0727 : integer;
		variable a0728 : integer;
		variable a0729 : integer;
		variable a0730 : integer;
		variable a0731 : integer;
		variable a0732 : integer;
		variable a0733 : integer;
		variable a0734 : integer;
		variable a0735 : integer;
		variable a0736 : integer;
		variable a0737 : integer;
		variable a0738 : integer;
		variable a0739 : integer;
		variable a0740 : integer;
		variable a0741 : integer;
		variable a0742 : integer;
		variable a0743 : integer;
		variable a0744 : integer;
		variable a0745 : integer;
		variable a0746 : integer;
		variable a0747 : integer;
		variable a0748 : integer;
		variable a0749 : integer;
		variable a0750 : integer;
		variable a0751 : integer;
		variable a0752 : integer;
		variable a0753 : integer;
		variable a0754 : integer;
		variable a0755 : integer;
		variable a0756 : integer;
		variable a0757 : integer;
		variable a0758 : integer;
		variable a0759 : integer;
		variable a0760 : integer;
		variable a0761 : integer;
		variable a0762 : integer;
		variable a0763 : integer;
		variable a0764 : integer;
		variable a0765 : integer;
		variable a0766 : integer;
		variable a0767 : integer;
		variable a0768 : integer;
		variable a0769 : integer;
		variable a0770 : integer;
		variable a0771 : integer;
		variable a0772 : integer;
		variable a0773 : integer;
		variable a0774 : integer;
		variable a0775 : integer;
		variable a0776 : integer;
		variable a0777 : integer;
		variable a0778 : integer;
		variable a0779 : integer;
		variable a0780 : integer;
		variable a0781 : integer;
		variable a0782 : integer;
		variable a0783 : integer;
		variable a0784 : integer;
		variable a0785 : integer;
		variable a0786 : integer;
		variable a0787 : integer;
		variable a0788 : integer;
		variable a0789 : integer;
		variable a0790 : integer;
		variable a0791 : integer;
		variable a0792 : integer;
		variable a0793 : integer;
		variable a0794 : integer;
		variable a0795 : integer;
		variable a0796 : integer;
		variable a0797 : integer;
		variable a0798 : integer;
		variable a0799 : integer;
		variable a0800 : integer;
		variable a0801 : integer;
		variable a0802 : integer;
		variable a0803 : integer;
		variable a0804 : integer;
		variable a0805 : integer;
		variable a0806 : integer;
		variable a0807 : integer;
		variable a0808 : integer;
		variable a0809 : integer;
		variable a0810 : integer;
		variable a0811 : integer;
		variable a0812 : integer;
		variable a0813 : integer;
		variable a0814 : integer;
		variable a0815 : integer;
		variable a0816 : integer;
		variable a0817 : integer;
		variable a0818 : integer;
		variable a0819 : integer;
		variable a0820 : integer;
		variable a0821 : integer;
		variable a0822 : integer;
		variable a0823 : integer;
		variable a0824 : integer;
		variable a0825 : integer;
		variable a0826 : integer;
		variable a0827 : integer;
		variable a0828 : integer;
		variable a0829 : integer;
		variable a0830 : integer;
		variable a0831 : integer;
		variable a0832 : integer;
		variable a0833 : integer;
		variable a0834 : integer;
		variable a0835 : integer;
		variable a0836 : integer;
		variable a0837 : integer;
		variable a0838 : integer;
		variable a0839 : integer;
		variable a0840 : integer;
		variable a0841 : integer;
		variable a0842 : integer;
		variable a0843 : integer;
		variable a0844 : integer;
		variable a0845 : integer;
		variable a0846 : integer;
		variable a0847 : integer;
		variable a0848 : integer;
		variable a0849 : integer;
		variable a0850 : integer;
		variable a0851 : integer;
		variable a0852 : integer;
		variable a0853 : integer;
		variable a0854 : integer;
		variable a0855 : integer;
		variable a0856 : integer;
		variable a0857 : integer;
		variable a0858 : integer;
		variable a0859 : integer;
		variable a0860 : integer;
		variable a0861 : integer;
		variable a0862 : integer;
		variable a0863 : integer;
		variable a0864 : integer;
		variable a0865 : integer;
		variable a0866 : integer;
		variable a0867 : integer;
		variable a0868 : integer;
		variable a0869 : integer;
		variable a0870 : integer;
		variable a0871 : integer;
		variable a0872 : integer;
		variable a0873 : integer;
		variable a0874 : integer;
		variable a0875 : integer;
		variable a0876 : integer;
		variable a0877 : integer;
		variable a0878 : integer;
		variable a0879 : integer;
		variable a0880 : integer;
		variable a0881 : integer;
		variable a0882 : integer;
		variable a0883 : integer;
		variable a0884 : integer;
		variable a0885 : integer;
		variable a0886 : integer;
		variable a0887 : integer;
		variable a0888 : integer;
		variable a0889 : integer;
		variable a0890 : integer;
		variable a0891 : integer;
		variable a0892 : integer;
		variable a0893 : integer;
		variable a0894 : integer;
		variable a0895 : integer;
		variable a0896 : integer;
		variable a0897 : integer;
		variable a0898 : integer;
		variable a0899 : integer;
		variable a0900 : integer;
		variable a0901 : integer;
		variable a0902 : integer;
		variable a0903 : integer;
		variable a0904 : integer;
		variable a0905 : integer;
		variable a0906 : integer;
		variable a0907 : integer;
		variable a0908 : integer;
		variable a0909 : integer;
		variable a0910 : integer;
		variable a0911 : integer;
		variable a0912 : integer;
		variable a0913 : integer;
		variable a0914 : integer;
		variable a0915 : integer;
		variable a0916 : integer;
		variable a0917 : integer;
		variable a0918 : integer;
		variable a0919 : integer;
		variable a0920 : integer;
		variable a0921 : integer;
		variable a0922 : integer;
		variable a0923 : integer;
		variable a0924 : integer;
		variable a0925 : integer;
		variable a0926 : integer;
		variable a0927 : integer;
		variable a0928 : integer;
		variable a0929 : integer;
		variable a0930 : integer;
		variable a0931 : integer;
		variable a0932 : integer;
		variable a0933 : integer;
		variable a0934 : integer;
		variable a0935 : integer;
		variable a0936 : integer;
		variable a0937 : integer;
		variable a0938 : integer;
		variable a0939 : integer;
		variable a0940 : integer;
		variable a0941 : integer;
		variable a0942 : integer;
		variable a0943 : integer;
		variable a0944 : integer;
		variable a0945 : integer;
		variable a0946 : integer;
		variable a0947 : integer;
		variable a0948 : integer;
		variable a0949 : integer;
		variable a0950 : integer;
		variable a0951 : integer;
		variable a0952 : integer;
		variable a0953 : integer;
		variable a0954 : integer;
		variable a0955 : integer;
		variable a0956 : integer;
		variable a0957 : integer;
		variable a0958 : integer;
		variable a0959 : integer;
		variable a0960 : integer;
		variable a0961 : integer;
		variable a0962 : integer;
		variable a0963 : integer;
		variable a0964 : integer;
		variable a0965 : integer;
		variable a0966 : integer;
		variable a0967 : integer;
		variable a0968 : integer;
		variable a0969 : integer;
		variable a0970 : integer;
		variable a0971 : integer;
		variable a0972 : integer;
		variable a0973 : integer;
		variable a0974 : integer;
		variable a0975 : integer;
		variable a0976 : integer;
		variable a0977 : integer;
		variable a0978 : integer;
		variable a0979 : integer;
		variable a0980 : integer;
		variable a0981 : integer;
		variable a0982 : integer;
		variable a0983 : integer;
		variable a0984 : integer;
		variable a0985 : integer;
		variable a0986 : integer;
		variable a0987 : integer;
		variable a0988 : integer;
		variable a0989 : integer;
		variable a0990 : integer;
		variable a0991 : integer;
		variable a0992 : integer;
		variable a0993 : integer;
		variable a0994 : integer;
		variable a0995 : integer;
		variable a0996 : integer;
		variable a0997 : integer;
		variable a0998 : integer;
		variable a0999 : integer;
		variable a1000 : integer;
	begin
		a0502 := clk;
		a0503 := clk;
		a0504 := clk;
		a0505 := clk;
		a0506 := clk;
		a0507 := clk;
		a0508 := clk;
		a0509 := clk;
		a0510 := clk;
		a0511 := clk;
		a0512 := clk;
		a0513 := clk;
		a0514 := clk;
		a0515 := clk;
		a0516 := clk;
		a0517 := clk;
		a0518 := clk;
		a0519 := clk;
		a0520 := clk;
		a0521 := clk;
		a0522 := clk;
		a0523 := clk;
		a0524 := clk;
		a0525 := clk;
		a0526 := clk;
		a0527 := clk;
		a0528 := clk;
		a0529 := clk;
		a0530 := clk;
		a0531 := clk;
		a0532 := clk;
		a0533 := clk;
		a0534 := clk;
		a0535 := clk;
		a0536 := clk;
		a0537 := clk;
		a0538 := clk;
		a0539 := clk;
		a0540 := clk;
		a0541 := clk;
		a0542 := clk;
		a0543 := clk;
		a0544 := clk;
		a0545 := clk;
		a0546 := clk;
		a0547 := clk;
		a0548 := clk;
		a0549 := clk;
		a0550 := clk;
		a0551 := clk;
		a0552 := clk;
		a0553 := clk;
		a0554 := clk;
		a0555 := clk;
		a0556 := clk;
		a0557 := clk;
		a0558 := clk;
		a0559 := clk;
		a0560 := clk;
		a0561 := clk;
		a0562 := clk;
		a0563 := clk;
		a0564 := clk;
		a0565 := clk;
		a0566 := clk;
		a0567 := clk;
		a0568 := clk;
		a0569 := clk;
		a0570 := clk;
		a0571 := clk;
		a0572 := clk;
		a0573 := clk;
		a0574 := clk;
		a0575 := clk;
		a0576 := clk;
		a0577 := clk;
		a0578 := clk;
		a0579 := clk;
		a0580 := clk;
		a0581 := clk;
		a0582 := clk;
		a0583 := clk;
		a0584 := clk;
		a0585 := clk;
		a0586 := clk;
		a0587 := clk;
		a0588 := clk;
		a0589 := clk;
		a0590 := clk;
		a0591 := clk;
		a0592 := clk;
		a0593 := clk;
		a0594 := clk;
		a0595 := clk;
		a0596 := clk;
		a0597 := clk;
		a0598 := clk;
		a0599 := clk;
		a0600 := clk;
		a0601 := clk;
		a0602 := clk;
		a0603 := clk;
		a0604 := clk;
		a0605 := clk;
		a0606 := clk;
		a0607 := clk;
		a0608 := clk;
		a0609 := clk;
		a0610 := clk;
		a0611 := clk;
		a0612 := clk;
		a0613 := clk;
		a0614 := clk;
		a0615 := clk;
		a0616 := clk;
		a0617 := clk;
		a0618 := clk;
		a0619 := clk;
		a0620 := clk;
		a0621 := clk;
		a0622 := clk;
		a0623 := clk;
		a0624 := clk;
		a0625 := clk;
		a0626 := clk;
		a0627 := clk;
		a0628 := clk;
		a0629 := clk;
		a0630 := clk;
		a0631 := clk;
		a0632 := clk;
		a0633 := clk;
		a0634 := clk;
		a0635 := clk;
		a0636 := clk;
		a0637 := clk;
		a0638 := clk;
		a0639 := clk;
		a0640 := clk;
		a0641 := clk;
		a0642 := clk;
		a0643 := clk;
		a0644 := clk;
		a0645 := clk;
		a0646 := clk;
		a0647 := clk;
		a0648 := clk;
		a0649 := clk;
		a0650 := clk;
		a0651 := clk;
		a0652 := clk;
		a0653 := clk;
		a0654 := clk;
		a0655 := clk;
		a0656 := clk;
		a0657 := clk;
		a0658 := clk;
		a0659 := clk;
		a0660 := clk;
		a0661 := clk;
		a0662 := clk;
		a0663 := clk;
		a0664 := clk;
		a0665 := clk;
		a0666 := clk;
		a0667 := clk;
		a0668 := clk;
		a0669 := clk;
		a0670 := clk;
		a0671 := clk;
		a0672 := clk;
		a0673 := clk;
		a0674 := clk;
		a0675 := clk;
		a0676 := clk;
		a0677 := clk;
		a0678 := clk;
		a0679 := clk;
		a0680 := clk;
		a0681 := clk;
		a0682 := clk;
		a0683 := clk;
		a0684 := clk;
		a0685 := clk;
		a0686 := clk;
		a0687 := clk;
		a0688 := clk;
		a0689 := clk;
		a0690 := clk;
		a0691 := clk;
		a0692 := clk;
		a0693 := clk;
		a0694 := clk;
		a0695 := clk;
		a0696 := clk;
		a0697 := clk;
		a0698 := clk;
		a0699 := clk;
		a0700 := clk;
		a0701 := clk;
		a0702 := clk;
		a0703 := clk;
		a0704 := clk;
		a0705 := clk;
		a0706 := clk;
		a0707 := clk;
		a0708 := clk;
		a0709 := clk;
		a0710 := clk;
		a0711 := clk;
		a0712 := clk;
		a0713 := clk;
		a0714 := clk;
		a0715 := clk;
		a0716 := clk;
		a0717 := clk;
		a0718 := clk;
		a0719 := clk;
		a0720 := clk;
		a0721 := clk;
		a0722 := clk;
		a0723 := clk;
		a0724 := clk;
		a0725 := clk;
		a0726 := clk;
		a0727 := clk;
		a0728 := clk;
		a0729 := clk;
		a0730 := clk;
		a0731 := clk;
		a0732 := clk;
		a0733 := clk;
		a0734 := clk;
		a0735 := clk;
		a0736 := clk;
		a0737 := clk;
		a0738 := clk;
		a0739 := clk;
		a0740 := clk;
		a0741 := clk;
		a0742 := clk;
		a0743 := clk;
		a0744 := clk;
		a0745 := clk;
		a0746 := clk;
		a0747 := clk;
		a0748 := clk;
		a0749 := clk;
		a0750 := clk;
		a0751 := clk;
		a0752 := clk;
		a0753 := clk;
		a0754 := clk;
		a0755 := clk;
		a0756 := clk;
		a0757 := clk;
		a0758 := clk;
		a0759 := clk;
		a0760 := clk;
		a0761 := clk;
		a0762 := clk;
		a0763 := clk;
		a0764 := clk;
		a0765 := clk;
		a0766 := clk;
		a0767 := clk;
		a0768 := clk;
		a0769 := clk;
		a0770 := clk;
		a0771 := clk;
		a0772 := clk;
		a0773 := clk;
		a0774 := clk;
		a0775 := clk;
		a0776 := clk;
		a0777 := clk;
		a0778 := clk;
		a0779 := clk;
		a0780 := clk;
		a0781 := clk;
		a0782 := clk;
		a0783 := clk;
		a0784 := clk;
		a0785 := clk;
		a0786 := clk;
		a0787 := clk;
		a0788 := clk;
		a0789 := clk;
		a0790 := clk;
		a0791 := clk;
		a0792 := clk;
		a0793 := clk;
		a0794 := clk;
		a0795 := clk;
		a0796 := clk;
		a0797 := clk;
		a0798 := clk;
		a0799 := clk;
		a0800 := clk;
		a0801 := clk;
		a0802 := clk;
		a0803 := clk;
		a0804 := clk;
		a0805 := clk;
		a0806 := clk;
		a0807 := clk;
		a0808 := clk;
		a0809 := clk;
		a0810 := clk;
		a0811 := clk;
		a0812 := clk;
		a0813 := clk;
		a0814 := clk;
		a0815 := clk;
		a0816 := clk;
		a0817 := clk;
		a0818 := clk;
		a0819 := clk;
		a0820 := clk;
		a0821 := clk;
		a0822 := clk;
		a0823 := clk;
		a0824 := clk;
		a0825 := clk;
		a0826 := clk;
		a0827 := clk;
		a0828 := clk;
		a0829 := clk;
		a0830 := clk;
		a0831 := clk;
		a0832 := clk;
		a0833 := clk;
		a0834 := clk;
		a0835 := clk;
		a0836 := clk;
		a0837 := clk;
		a0838 := clk;
		a0839 := clk;
		a0840 := clk;
		a0841 := clk;
		a0842 := clk;
		a0843 := clk;
		a0844 := clk;
		a0845 := clk;
		a0846 := clk;
		a0847 := clk;
		a0848 := clk;
		a0849 := clk;
		a0850 := clk;
		a0851 := clk;
		a0852 := clk;
		a0853 := clk;
		a0854 := clk;
		a0855 := clk;
		a0856 := clk;
		a0857 := clk;
		a0858 := clk;
		a0859 := clk;
		a0860 := clk;
		a0861 := clk;
		a0862 := clk;
		a0863 := clk;
		a0864 := clk;
		a0865 := clk;
		a0866 := clk;
		a0867 := clk;
		a0868 := clk;
		a0869 := clk;
		a0870 := clk;
		a0871 := clk;
		a0872 := clk;
		a0873 := clk;
		a0874 := clk;
		a0875 := clk;
		a0876 := clk;
		a0877 := clk;
		a0878 := clk;
		a0879 := clk;
		a0880 := clk;
		a0881 := clk;
		a0882 := clk;
		a0883 := clk;
		a0884 := clk;
		a0885 := clk;
		a0886 := clk;
		a0887 := clk;
		a0888 := clk;
		a0889 := clk;
		a0890 := clk;
		a0891 := clk;
		a0892 := clk;
		a0893 := clk;
		a0894 := clk;
		a0895 := clk;
		a0896 := clk;
		a0897 := clk;
		a0898 := clk;
		a0899 := clk;
		a0900 := clk;
		a0901 := clk;
		a0902 := clk;
		a0903 := clk;
		a0904 := clk;
		a0905 := clk;
		a0906 := clk;
		a0907 := clk;
		a0908 := clk;
		a0909 := clk;
		a0910 := clk;
		a0911 := clk;
		a0912 := clk;
		a0913 := clk;
		a0914 := clk;
		a0915 := clk;
		a0916 := clk;
		a0917 := clk;
		a0918 := clk;
		a0919 := clk;
		a0920 := clk;
		a0921 := clk;
		a0922 := clk;
		a0923 := clk;
		a0924 := clk;
		a0925 := clk;
		a0926 := clk;
		a0927 := clk;
		a0928 := clk;
		a0929 := clk;
		a0930 := clk;
		a0931 := clk;
		a0932 := clk;
		a0933 := clk;
		a0934 := clk;
		a0935 := clk;
		a0936 := clk;
		a0937 := clk;
		a0938 := clk;
		a0939 := clk;
		a0940 := clk;
		a0941 := clk;
		a0942 := clk;
		a0943 := clk;
		a0944 := clk;
		a0945 := clk;
		a0946 := clk;
		a0947 := clk;
		a0948 := clk;
		a0949 := clk;
		a0950 := clk;
		a0951 := clk;
		a0952 := clk;
		a0953 := clk;
		a0954 := clk;
		a0955 := clk;
		a0956 := clk;
		a0957 := clk;
		a0958 := clk;
		a0959 := clk;
		a0960 := clk;
		a0961 := clk;
		a0962 := clk;
		a0963 := clk;
		a0964 := clk;
		a0965 := clk;
		a0966 := clk;
		a0967 := clk;
		a0968 := clk;
		a0969 := clk;
		a0970 := clk;
		a0971 := clk;
		a0972 := clk;
		a0973 := clk;
		a0974 := clk;
		a0975 := clk;
		a0976 := clk;
		a0977 := clk;
		a0978 := clk;
		a0979 := clk;
		a0980 := clk;
		a0981 := clk;
		a0982 := clk;
		a0983 := clk;
		a0984 := clk;
		a0985 := clk;
		a0986 := clk;
		a0987 := clk;
		a0988 := clk;
		a0989 := clk;
		a0990 := clk;
		a0991 := clk;
		a0992 := clk;
		a0993 := clk;
		a0994 := clk;
		a0995 := clk;
		a0996 := clk;
		a0997 := clk;
		a0998 := clk;
		a0999 := clk;
		a1000 := clk;
	--}}}
	end process;

	main1: process(clk)
		--{{{
		variable a0502 : integer;
		variable a0503 : integer;
		variable a0504 : integer;
		variable a0505 : integer;
		variable a0506 : integer;
		variable a0507 : integer;
		variable a0508 : integer;
		variable a0509 : integer;
		variable a0510 : integer;
		variable a0511 : integer;
		variable a0512 : integer;
		variable a0513 : integer;
		variable a0514 : integer;
		variable a0515 : integer;
		variable a0516 : integer;
		variable a0517 : integer;
		variable a0518 : integer;
		variable a0519 : integer;
		variable a0520 : integer;
		variable a0521 : integer;
		variable a0522 : integer;
		variable a0523 : integer;
		variable a0524 : integer;
		variable a0525 : integer;
		variable a0526 : integer;
		variable a0527 : integer;
		variable a0528 : integer;
		variable a0529 : integer;
		variable a0530 : integer;
		variable a0531 : integer;
		variable a0532 : integer;
		variable a0533 : integer;
		variable a0534 : integer;
		variable a0535 : integer;
		variable a0536 : integer;
		variable a0537 : integer;
		variable a0538 : integer;
		variable a0539 : integer;
		variable a0540 : integer;
		variable a0541 : integer;
		variable a0542 : integer;
		variable a0543 : integer;
		variable a0544 : integer;
		variable a0545 : integer;
		variable a0546 : integer;
		variable a0547 : integer;
		variable a0548 : integer;
		variable a0549 : integer;
		variable a0550 : integer;
		variable a0551 : integer;
		variable a0552 : integer;
		variable a0553 : integer;
		variable a0554 : integer;
		variable a0555 : integer;
		variable a0556 : integer;
		variable a0557 : integer;
		variable a0558 : integer;
		variable a0559 : integer;
		variable a0560 : integer;
		variable a0561 : integer;
		variable a0562 : integer;
		variable a0563 : integer;
		variable a0564 : integer;
		variable a0565 : integer;
		variable a0566 : integer;
		variable a0567 : integer;
		variable a0568 : integer;
		variable a0569 : integer;
		variable a0570 : integer;
		variable a0571 : integer;
		variable a0572 : integer;
		variable a0573 : integer;
		variable a0574 : integer;
		variable a0575 : integer;
		variable a0576 : integer;
		variable a0577 : integer;
		variable a0578 : integer;
		variable a0579 : integer;
		variable a0580 : integer;
		variable a0581 : integer;
		variable a0582 : integer;
		variable a0583 : integer;
		variable a0584 : integer;
		variable a0585 : integer;
		variable a0586 : integer;
		variable a0587 : integer;
		variable a0588 : integer;
		variable a0589 : integer;
		variable a0590 : integer;
		variable a0591 : integer;
		variable a0592 : integer;
		variable a0593 : integer;
		variable a0594 : integer;
		variable a0595 : integer;
		variable a0596 : integer;
		variable a0597 : integer;
		variable a0598 : integer;
		variable a0599 : integer;
		variable a0600 : integer;
		variable a0601 : integer;
		variable a0602 : integer;
		variable a0603 : integer;
		variable a0604 : integer;
		variable a0605 : integer;
		variable a0606 : integer;
		variable a0607 : integer;
		variable a0608 : integer;
		variable a0609 : integer;
		variable a0610 : integer;
		variable a0611 : integer;
		variable a0612 : integer;
		variable a0613 : integer;
		variable a0614 : integer;
		variable a0615 : integer;
		variable a0616 : integer;
		variable a0617 : integer;
		variable a0618 : integer;
		variable a0619 : integer;
		variable a0620 : integer;
		variable a0621 : integer;
		variable a0622 : integer;
		variable a0623 : integer;
		variable a0624 : integer;
		variable a0625 : integer;
		variable a0626 : integer;
		variable a0627 : integer;
		variable a0628 : integer;
		variable a0629 : integer;
		variable a0630 : integer;
		variable a0631 : integer;
		variable a0632 : integer;
		variable a0633 : integer;
		variable a0634 : integer;
		variable a0635 : integer;
		variable a0636 : integer;
		variable a0637 : integer;
		variable a0638 : integer;
		variable a0639 : integer;
		variable a0640 : integer;
		variable a0641 : integer;
		variable a0642 : integer;
		variable a0643 : integer;
		variable a0644 : integer;
		variable a0645 : integer;
		variable a0646 : integer;
		variable a0647 : integer;
		variable a0648 : integer;
		variable a0649 : integer;
		variable a0650 : integer;
		variable a0651 : integer;
		variable a0652 : integer;
		variable a0653 : integer;
		variable a0654 : integer;
		variable a0655 : integer;
		variable a0656 : integer;
		variable a0657 : integer;
		variable a0658 : integer;
		variable a0659 : integer;
		variable a0660 : integer;
		variable a0661 : integer;
		variable a0662 : integer;
		variable a0663 : integer;
		variable a0664 : integer;
		variable a0665 : integer;
		variable a0666 : integer;
		variable a0667 : integer;
		variable a0668 : integer;
		variable a0669 : integer;
		variable a0670 : integer;
		variable a0671 : integer;
		variable a0672 : integer;
		variable a0673 : integer;
		variable a0674 : integer;
		variable a0675 : integer;
		variable a0676 : integer;
		variable a0677 : integer;
		variable a0678 : integer;
		variable a0679 : integer;
		variable a0680 : integer;
		variable a0681 : integer;
		variable a0682 : integer;
		variable a0683 : integer;
		variable a0684 : integer;
		variable a0685 : integer;
		variable a0686 : integer;
		variable a0687 : integer;
		variable a0688 : integer;
		variable a0689 : integer;
		variable a0690 : integer;
		variable a0691 : integer;
		variable a0692 : integer;
		variable a0693 : integer;
		variable a0694 : integer;
		variable a0695 : integer;
		variable a0696 : integer;
		variable a0697 : integer;
		variable a0698 : integer;
		variable a0699 : integer;
		variable a0700 : integer;
		variable a0701 : integer;
		variable a0702 : integer;
		variable a0703 : integer;
		variable a0704 : integer;
		variable a0705 : integer;
		variable a0706 : integer;
		variable a0707 : integer;
		variable a0708 : integer;
		variable a0709 : integer;
		variable a0710 : integer;
		variable a0711 : integer;
		variable a0712 : integer;
		variable a0713 : integer;
		variable a0714 : integer;
		variable a0715 : integer;
		variable a0716 : integer;
		variable a0717 : integer;
		variable a0718 : integer;
		variable a0719 : integer;
		variable a0720 : integer;
		variable a0721 : integer;
		variable a0722 : integer;
		variable a0723 : integer;
		variable a0724 : integer;
		variable a0725 : integer;
		variable a0726 : integer;
		variable a0727 : integer;
		variable a0728 : integer;
		variable a0729 : integer;
		variable a0730 : integer;
		variable a0731 : integer;
		variable a0732 : integer;
		variable a0733 : integer;
		variable a0734 : integer;
		variable a0735 : integer;
		variable a0736 : integer;
		variable a0737 : integer;
		variable a0738 : integer;
		variable a0739 : integer;
		variable a0740 : integer;
		variable a0741 : integer;
		variable a0742 : integer;
		variable a0743 : integer;
		variable a0744 : integer;
		variable a0745 : integer;
		variable a0746 : integer;
		variable a0747 : integer;
		variable a0748 : integer;
		variable a0749 : integer;
		variable a0750 : integer;
		variable a0751 : integer;
		variable a0752 : integer;
		variable a0753 : integer;
		variable a0754 : integer;
		variable a0755 : integer;
		variable a0756 : integer;
		variable a0757 : integer;
		variable a0758 : integer;
		variable a0759 : integer;
		variable a0760 : integer;
		variable a0761 : integer;
		variable a0762 : integer;
		variable a0763 : integer;
		variable a0764 : integer;
		variable a0765 : integer;
		variable a0766 : integer;
		variable a0767 : integer;
		variable a0768 : integer;
		variable a0769 : integer;
		variable a0770 : integer;
		variable a0771 : integer;
		variable a0772 : integer;
		variable a0773 : integer;
		variable a0774 : integer;
		variable a0775 : integer;
		variable a0776 : integer;
		variable a0777 : integer;
		variable a0778 : integer;
		variable a0779 : integer;
		variable a0780 : integer;
		variable a0781 : integer;
		variable a0782 : integer;
		variable a0783 : integer;
		variable a0784 : integer;
		variable a0785 : integer;
		variable a0786 : integer;
		variable a0787 : integer;
		variable a0788 : integer;
		variable a0789 : integer;
		variable a0790 : integer;
		variable a0791 : integer;
		variable a0792 : integer;
		variable a0793 : integer;
		variable a0794 : integer;
		variable a0795 : integer;
		variable a0796 : integer;
		variable a0797 : integer;
		variable a0798 : integer;
		variable a0799 : integer;
		variable a0800 : integer;
		variable a0801 : integer;
		variable a0802 : integer;
		variable a0803 : integer;
		variable a0804 : integer;
		variable a0805 : integer;
		variable a0806 : integer;
		variable a0807 : integer;
		variable a0808 : integer;
		variable a0809 : integer;
		variable a0810 : integer;
		variable a0811 : integer;
		variable a0812 : integer;
		variable a0813 : integer;
		variable a0814 : integer;
		variable a0815 : integer;
		variable a0816 : integer;
		variable a0817 : integer;
		variable a0818 : integer;
		variable a0819 : integer;
		variable a0820 : integer;
		variable a0821 : integer;
		variable a0822 : integer;
		variable a0823 : integer;
		variable a0824 : integer;
		variable a0825 : integer;
		variable a0826 : integer;
		variable a0827 : integer;
		variable a0828 : integer;
		variable a0829 : integer;
		variable a0830 : integer;
		variable a0831 : integer;
		variable a0832 : integer;
		variable a0833 : integer;
		variable a0834 : integer;
		variable a0835 : integer;
		variable a0836 : integer;
		variable a0837 : integer;
		variable a0838 : integer;
		variable a0839 : integer;
		variable a0840 : integer;
		variable a0841 : integer;
		variable a0842 : integer;
		variable a0843 : integer;
		variable a0844 : integer;
		variable a0845 : integer;
		variable a0846 : integer;
		variable a0847 : integer;
		variable a0848 : integer;
		variable a0849 : integer;
		variable a0850 : integer;
		variable a0851 : integer;
		variable a0852 : integer;
		variable a0853 : integer;
		variable a0854 : integer;
		variable a0855 : integer;
		variable a0856 : integer;
		variable a0857 : integer;
		variable a0858 : integer;
		variable a0859 : integer;
		variable a0860 : integer;
		variable a0861 : integer;
		variable a0862 : integer;
		variable a0863 : integer;
		variable a0864 : integer;
		variable a0865 : integer;
		variable a0866 : integer;
		variable a0867 : integer;
		variable a0868 : integer;
		variable a0869 : integer;
		variable a0870 : integer;
		variable a0871 : integer;
		variable a0872 : integer;
		variable a0873 : integer;
		variable a0874 : integer;
		variable a0875 : integer;
		variable a0876 : integer;
		variable a0877 : integer;
		variable a0878 : integer;
		variable a0879 : integer;
		variable a0880 : integer;
		variable a0881 : integer;
		variable a0882 : integer;
		variable a0883 : integer;
		variable a0884 : integer;
		variable a0885 : integer;
		variable a0886 : integer;
		variable a0887 : integer;
		variable a0888 : integer;
		variable a0889 : integer;
		variable a0890 : integer;
		variable a0891 : integer;
		variable a0892 : integer;
		variable a0893 : integer;
		variable a0894 : integer;
		variable a0895 : integer;
		variable a0896 : integer;
		variable a0897 : integer;
		variable a0898 : integer;
		variable a0899 : integer;
		variable a0900 : integer;
		variable a0901 : integer;
		variable a0902 : integer;
		variable a0903 : integer;
		variable a0904 : integer;
		variable a0905 : integer;
		variable a0906 : integer;
		variable a0907 : integer;
		variable a0908 : integer;
		variable a0909 : integer;
		variable a0910 : integer;
		variable a0911 : integer;
		variable a0912 : integer;
		variable a0913 : integer;
		variable a0914 : integer;
		variable a0915 : integer;
		variable a0916 : integer;
		variable a0917 : integer;
		variable a0918 : integer;
		variable a0919 : integer;
		variable a0920 : integer;
		variable a0921 : integer;
		variable a0922 : integer;
		variable a0923 : integer;
		variable a0924 : integer;
		variable a0925 : integer;
		variable a0926 : integer;
		variable a0927 : integer;
		variable a0928 : integer;
		variable a0929 : integer;
		variable a0930 : integer;
		variable a0931 : integer;
		variable a0932 : integer;
		variable a0933 : integer;
		variable a0934 : integer;
		variable a0935 : integer;
		variable a0936 : integer;
		variable a0937 : integer;
		variable a0938 : integer;
		variable a0939 : integer;
		variable a0940 : integer;
		variable a0941 : integer;
		variable a0942 : integer;
		variable a0943 : integer;
		variable a0944 : integer;
		variable a0945 : integer;
		variable a0946 : integer;
		variable a0947 : integer;
		variable a0948 : integer;
		variable a0949 : integer;
		variable a0950 : integer;
		variable a0951 : integer;
		variable a0952 : integer;
		variable a0953 : integer;
		variable a0954 : integer;
		variable a0955 : integer;
		variable a0956 : integer;
		variable a0957 : integer;
		variable a0958 : integer;
		variable a0959 : integer;
		variable a0960 : integer;
		variable a0961 : integer;
		variable a0962 : integer;
		variable a0963 : integer;
		variable a0964 : integer;
		variable a0965 : integer;
		variable a0966 : integer;
		variable a0967 : integer;
		variable a0968 : integer;
		variable a0969 : integer;
		variable a0970 : integer;
		variable a0971 : integer;
		variable a0972 : integer;
		variable a0973 : integer;
		variable a0974 : integer;
		variable a0975 : integer;
		variable a0976 : integer;
		variable a0977 : integer;
		variable a0978 : integer;
		variable a0979 : integer;
		variable a0980 : integer;
		variable a0981 : integer;
		variable a0982 : integer;
		variable a0983 : integer;
		variable a0984 : integer;
		variable a0985 : integer;
		variable a0986 : integer;
		variable a0987 : integer;
		variable a0988 : integer;
		variable a0989 : integer;
		variable a0990 : integer;
		variable a0991 : integer;
		variable a0992 : integer;
		variable a0993 : integer;
		variable a0994 : integer;
		variable a0995 : integer;
		variable a0996 : integer;
		variable a0997 : integer;
		variable a0998 : integer;
		variable a0999 : integer;
		variable a1000 : integer;
	begin
		a0502 := clk;
		a0503 := clk;
		a0504 := clk;
		a0505 := clk;
		a0506 := clk;
		a0507 := clk;
		a0508 := clk;
		a0509 := clk;
		a0510 := clk;
		a0511 := clk;
		a0512 := clk;
		a0513 := clk;
		a0514 := clk;
		a0515 := clk;
		a0516 := clk;
		a0517 := clk;
		a0518 := clk;
		a0519 := clk;
		a0520 := clk;
		a0521 := clk;
		a0522 := clk;
		a0523 := clk;
		a0524 := clk;
		a0525 := clk;
		a0526 := clk;
		a0527 := clk;
		a0528 := clk;
		a0529 := clk;
		a0530 := clk;
		a0531 := clk;
		a0532 := clk;
		a0533 := clk;
		a0534 := clk;
		a0535 := clk;
		a0536 := clk;
		a0537 := clk;
		a0538 := clk;
		a0539 := clk;
		a0540 := clk;
		a0541 := clk;
		a0542 := clk;
		a0543 := clk;
		a0544 := clk;
		a0545 := clk;
		a0546 := clk;
		a0547 := clk;
		a0548 := clk;
		a0549 := clk;
		a0550 := clk;
		a0551 := clk;
		a0552 := clk;
		a0553 := clk;
		a0554 := clk;
		a0555 := clk;
		a0556 := clk;
		a0557 := clk;
		a0558 := clk;
		a0559 := clk;
		a0560 := clk;
		a0561 := clk;
		a0562 := clk;
		a0563 := clk;
		a0564 := clk;
		a0565 := clk;
		a0566 := clk;
		a0567 := clk;
		a0568 := clk;
		a0569 := clk;
		a0570 := clk;
		a0571 := clk;
		a0572 := clk;
		a0573 := clk;
		a0574 := clk;
		a0575 := clk;
		a0576 := clk;
		a0577 := clk;
		a0578 := clk;
		a0579 := clk;
		a0580 := clk;
		a0581 := clk;
		a0582 := clk;
		a0583 := clk;
		a0584 := clk;
		a0585 := clk;
		a0586 := clk;
		a0587 := clk;
		a0588 := clk;
		a0589 := clk;
		a0590 := clk;
		a0591 := clk;
		a0592 := clk;
		a0593 := clk;
		a0594 := clk;
		a0595 := clk;
		a0596 := clk;
		a0597 := clk;
		a0598 := clk;
		a0599 := clk;
		a0600 := clk;
		a0601 := clk;
		a0602 := clk;
		a0603 := clk;
		a0604 := clk;
		a0605 := clk;
		a0606 := clk;
		a0607 := clk;
		a0608 := clk;
		a0609 := clk;
		a0610 := clk;
		a0611 := clk;
		a0612 := clk;
		a0613 := clk;
		a0614 := clk;
		a0615 := clk;
		a0616 := clk;
		a0617 := clk;
		a0618 := clk;
		a0619 := clk;
		a0620 := clk;
		a0621 := clk;
		a0622 := clk;
		a0623 := clk;
		a0624 := clk;
		a0625 := clk;
		a0626 := clk;
		a0627 := clk;
		a0628 := clk;
		a0629 := clk;
		a0630 := clk;
		a0631 := clk;
		a0632 := clk;
		a0633 := clk;
		a0634 := clk;
		a0635 := clk;
		a0636 := clk;
		a0637 := clk;
		a0638 := clk;
		a0639 := clk;
		a0640 := clk;
		a0641 := clk;
		a0642 := clk;
		a0643 := clk;
		a0644 := clk;
		a0645 := clk;
		a0646 := clk;
		a0647 := clk;
		a0648 := clk;
		a0649 := clk;
		a0650 := clk;
		a0651 := clk;
		a0652 := clk;
		a0653 := clk;
		a0654 := clk;
		a0655 := clk;
		a0656 := clk;
		a0657 := clk;
		a0658 := clk;
		a0659 := clk;
		a0660 := clk;
		a0661 := clk;
		a0662 := clk;
		a0663 := clk;
		a0664 := clk;
		a0665 := clk;
		a0666 := clk;
		a0667 := clk;
		a0668 := clk;
		a0669 := clk;
		a0670 := clk;
		a0671 := clk;
		a0672 := clk;
		a0673 := clk;
		a0674 := clk;
		a0675 := clk;
		a0676 := clk;
		a0677 := clk;
		a0678 := clk;
		a0679 := clk;
		a0680 := clk;
		a0681 := clk;
		a0682 := clk;
		a0683 := clk;
		a0684 := clk;
		a0685 := clk;
		a0686 := clk;
		a0687 := clk;
		a0688 := clk;
		a0689 := clk;
		a0690 := clk;
		a0691 := clk;
		a0692 := clk;
		a0693 := clk;
		a0694 := clk;
		a0695 := clk;
		a0696 := clk;
		a0697 := clk;
		a0698 := clk;
		a0699 := clk;
		a0700 := clk;
		a0701 := clk;
		a0702 := clk;
		a0703 := clk;
		a0704 := clk;
		a0705 := clk;
		a0706 := clk;
		a0707 := clk;
		a0708 := clk;
		a0709 := clk;
		a0710 := clk;
		a0711 := clk;
		a0712 := clk;
		a0713 := clk;
		a0714 := clk;
		a0715 := clk;
		a0716 := clk;
		a0717 := clk;
		a0718 := clk;
		a0719 := clk;
		a0720 := clk;
		a0721 := clk;
		a0722 := clk;
		a0723 := clk;
		a0724 := clk;
		a0725 := clk;
		a0726 := clk;
		a0727 := clk;
		a0728 := clk;
		a0729 := clk;
		a0730 := clk;
		a0731 := clk;
		a0732 := clk;
		a0733 := clk;
		a0734 := clk;
		a0735 := clk;
		a0736 := clk;
		a0737 := clk;
		a0738 := clk;
		a0739 := clk;
		a0740 := clk;
		a0741 := clk;
		a0742 := clk;
		a0743 := clk;
		a0744 := clk;
		a0745 := clk;
		a0746 := clk;
		a0747 := clk;
		a0748 := clk;
		a0749 := clk;
		a0750 := clk;
		a0751 := clk;
		a0752 := clk;
		a0753 := clk;
		a0754 := clk;
		a0755 := clk;
		a0756 := clk;
		a0757 := clk;
		a0758 := clk;
		a0759 := clk;
		a0760 := clk;
		a0761 := clk;
		a0762 := clk;
		a0763 := clk;
		a0764 := clk;
		a0765 := clk;
		a0766 := clk;
		a0767 := clk;
		a0768 := clk;
		a0769 := clk;
		a0770 := clk;
		a0771 := clk;
		a0772 := clk;
		a0773 := clk;
		a0774 := clk;
		a0775 := clk;
		a0776 := clk;
		a0777 := clk;
		a0778 := clk;
		a0779 := clk;
		a0780 := clk;
		a0781 := clk;
		a0782 := clk;
		a0783 := clk;
		a0784 := clk;
		a0785 := clk;
		a0786 := clk;
		a0787 := clk;
		a0788 := clk;
		a0789 := clk;
		a0790 := clk;
		a0791 := clk;
		a0792 := clk;
		a0793 := clk;
		a0794 := clk;
		a0795 := clk;
		a0796 := clk;
		a0797 := clk;
		a0798 := clk;
		a0799 := clk;
		a0800 := clk;
		a0801 := clk;
		a0802 := clk;
		a0803 := clk;
		a0804 := clk;
		a0805 := clk;
		a0806 := clk;
		a0807 := clk;
		a0808 := clk;
		a0809 := clk;
		a0810 := clk;
		a0811 := clk;
		a0812 := clk;
		a0813 := clk;
		a0814 := clk;
		a0815 := clk;
		a0816 := clk;
		a0817 := clk;
		a0818 := clk;
		a0819 := clk;
		a0820 := clk;
		a0821 := clk;
		a0822 := clk;
		a0823 := clk;
		a0824 := clk;
		a0825 := clk;
		a0826 := clk;
		a0827 := clk;
		a0828 := clk;
		a0829 := clk;
		a0830 := clk;
		a0831 := clk;
		a0832 := clk;
		a0833 := clk;
		a0834 := clk;
		a0835 := clk;
		a0836 := clk;
		a0837 := clk;
		a0838 := clk;
		a0839 := clk;
		a0840 := clk;
		a0841 := clk;
		a0842 := clk;
		a0843 := clk;
		a0844 := clk;
		a0845 := clk;
		a0846 := clk;
		a0847 := clk;
		a0848 := clk;
		a0849 := clk;
		a0850 := clk;
		a0851 := clk;
		a0852 := clk;
		a0853 := clk;
		a0854 := clk;
		a0855 := clk;
		a0856 := clk;
		a0857 := clk;
		a0858 := clk;
		a0859 := clk;
		a0860 := clk;
		a0861 := clk;
		a0862 := clk;
		a0863 := clk;
		a0864 := clk;
		a0865 := clk;
		a0866 := clk;
		a0867 := clk;
		a0868 := clk;
		a0869 := clk;
		a0870 := clk;
		a0871 := clk;
		a0872 := clk;
		a0873 := clk;
		a0874 := clk;
		a0875 := clk;
		a0876 := clk;
		a0877 := clk;
		a0878 := clk;
		a0879 := clk;
		a0880 := clk;
		a0881 := clk;
		a0882 := clk;
		a0883 := clk;
		a0884 := clk;
		a0885 := clk;
		a0886 := clk;
		a0887 := clk;
		a0888 := clk;
		a0889 := clk;
		a0890 := clk;
		a0891 := clk;
		a0892 := clk;
		a0893 := clk;
		a0894 := clk;
		a0895 := clk;
		a0896 := clk;
		a0897 := clk;
		a0898 := clk;
		a0899 := clk;
		a0900 := clk;
		a0901 := clk;
		a0902 := clk;
		a0903 := clk;
		a0904 := clk;
		a0905 := clk;
		a0906 := clk;
		a0907 := clk;
		a0908 := clk;
		a0909 := clk;
		a0910 := clk;
		a0911 := clk;
		a0912 := clk;
		a0913 := clk;
		a0914 := clk;
		a0915 := clk;
		a0916 := clk;
		a0917 := clk;
		a0918 := clk;
		a0919 := clk;
		a0920 := clk;
		a0921 := clk;
		a0922 := clk;
		a0923 := clk;
		a0924 := clk;
		a0925 := clk;
		a0926 := clk;
		a0927 := clk;
		a0928 := clk;
		a0929 := clk;
		a0930 := clk;
		a0931 := clk;
		a0932 := clk;
		a0933 := clk;
		a0934 := clk;
		a0935 := clk;
		a0936 := clk;
		a0937 := clk;
		a0938 := clk;
		a0939 := clk;
		a0940 := clk;
		a0941 := clk;
		a0942 := clk;
		a0943 := clk;
		a0944 := clk;
		a0945 := clk;
		a0946 := clk;
		a0947 := clk;
		a0948 := clk;
		a0949 := clk;
		a0950 := clk;
		a0951 := clk;
		a0952 := clk;
		a0953 := clk;
		a0954 := clk;
		a0955 := clk;
		a0956 := clk;
		a0957 := clk;
		a0958 := clk;
		a0959 := clk;
		a0960 := clk;
		a0961 := clk;
		a0962 := clk;
		a0963 := clk;
		a0964 := clk;
		a0965 := clk;
		a0966 := clk;
		a0967 := clk;
		a0968 := clk;
		a0969 := clk;
		a0970 := clk;
		a0971 := clk;
		a0972 := clk;
		a0973 := clk;
		a0974 := clk;
		a0975 := clk;
		a0976 := clk;
		a0977 := clk;
		a0978 := clk;
		a0979 := clk;
		a0980 := clk;
		a0981 := clk;
		a0982 := clk;
		a0983 := clk;
		a0984 := clk;
		a0985 := clk;
		a0986 := clk;
		a0987 := clk;
		a0988 := clk;
		a0989 := clk;
		a0990 := clk;
		a0991 := clk;
		a0992 := clk;
		a0993 := clk;
		a0994 := clk;
		a0995 := clk;
		a0996 := clk;
		a0997 := clk;
		a0998 := clk;
		a0999 := clk;
		a1000 := clk;
	--}}}
	end process;

	terminator : process(clk)
	begin
		if clk >= CYCLES then
			assert false report "end of simulation" severity failure;
		-- else
		-- 	report "tick";
		end if;
	end process;

	clk <= (clk+1) after 1 us;
end;
