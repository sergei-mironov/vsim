entity ENT00001_Test_Bench is
end entity ENT00001_Test_Bench;

architecture arch of ENT00001_Test_Bench is
	signal clk : integer := 0;
	constant CYCLES : integer := 1000;
begin

	main: process(clk)
--{{{
		variable a0001 : integer;
		variable a0002 : integer;
		variable a0003 : integer;
		variable a0004 : integer;
		variable a0005 : integer;
		variable a0006 : integer;
		variable a0007 : integer;
		variable a0008 : integer;
		variable a0009 : integer;
		variable a0010 : integer;
		variable a0011 : integer;
		variable a0012 : integer;
		variable a0013 : integer;
		variable a0014 : integer;
		variable a0015 : integer;
		variable a0016 : integer;
		variable a0017 : integer;
		variable a0018 : integer;
		variable a0019 : integer;
		variable a0020 : integer;
		variable a0021 : integer;
		variable a0022 : integer;
		variable a0023 : integer;
		variable a0024 : integer;
		variable a0025 : integer;
		variable a0026 : integer;
		variable a0027 : integer;
		variable a0028 : integer;
		variable a0029 : integer;
		variable a0030 : integer;
		variable a0031 : integer;
		variable a0032 : integer;
		variable a0033 : integer;
		variable a0034 : integer;
		variable a0035 : integer;
		variable a0036 : integer;
		variable a0037 : integer;
		variable a0038 : integer;
		variable a0039 : integer;
		variable a0040 : integer;
		variable a0041 : integer;
		variable a0042 : integer;
		variable a0043 : integer;
		variable a0044 : integer;
		variable a0045 : integer;
		variable a0046 : integer;
		variable a0047 : integer;
		variable a0048 : integer;
		variable a0049 : integer;
		variable a0050 : integer;
		variable a0051 : integer;
		variable a0052 : integer;
		variable a0053 : integer;
		variable a0054 : integer;
		variable a0055 : integer;
		variable a0056 : integer;
		variable a0057 : integer;
		variable a0058 : integer;
		variable a0059 : integer;
		variable a0060 : integer;
		variable a0061 : integer;
		variable a0062 : integer;
		variable a0063 : integer;
		variable a0064 : integer;
		variable a0065 : integer;
		variable a0066 : integer;
		variable a0067 : integer;
		variable a0068 : integer;
		variable a0069 : integer;
		variable a0070 : integer;
		variable a0071 : integer;
		variable a0072 : integer;
		variable a0073 : integer;
		variable a0074 : integer;
		variable a0075 : integer;
		variable a0076 : integer;
		variable a0077 : integer;
		variable a0078 : integer;
		variable a0079 : integer;
		variable a0080 : integer;
		variable a0081 : integer;
		variable a0082 : integer;
		variable a0083 : integer;
		variable a0084 : integer;
		variable a0085 : integer;
		variable a0086 : integer;
		variable a0087 : integer;
		variable a0088 : integer;
		variable a0089 : integer;
		variable a0090 : integer;
		variable a0091 : integer;
		variable a0092 : integer;
		variable a0093 : integer;
		variable a0094 : integer;
		variable a0095 : integer;
		variable a0096 : integer;
		variable a0097 : integer;
		variable a0098 : integer;
		variable a0099 : integer;
		variable a0100 : integer;
		variable a0101 : integer;
		variable a0102 : integer;
		variable a0103 : integer;
		variable a0104 : integer;
		variable a0105 : integer;
		variable a0106 : integer;
		variable a0107 : integer;
		variable a0108 : integer;
		variable a0109 : integer;
		variable a0110 : integer;
		variable a0111 : integer;
		variable a0112 : integer;
		variable a0113 : integer;
		variable a0114 : integer;
		variable a0115 : integer;
		variable a0116 : integer;
		variable a0117 : integer;
		variable a0118 : integer;
		variable a0119 : integer;
		variable a0120 : integer;
		variable a0121 : integer;
		variable a0122 : integer;
		variable a0123 : integer;
		variable a0124 : integer;
		variable a0125 : integer;
		variable a0126 : integer;
		variable a0127 : integer;
		variable a0128 : integer;
		variable a0129 : integer;
		variable a0130 : integer;
		variable a0131 : integer;
		variable a0132 : integer;
		variable a0133 : integer;
		variable a0134 : integer;
		variable a0135 : integer;
		variable a0136 : integer;
		variable a0137 : integer;
		variable a0138 : integer;
		variable a0139 : integer;
		variable a0140 : integer;
		variable a0141 : integer;
		variable a0142 : integer;
		variable a0143 : integer;
		variable a0144 : integer;
		variable a0145 : integer;
		variable a0146 : integer;
		variable a0147 : integer;
		variable a0148 : integer;
		variable a0149 : integer;
		variable a0150 : integer;
		variable a0151 : integer;
		variable a0152 : integer;
		variable a0153 : integer;
		variable a0154 : integer;
		variable a0155 : integer;
		variable a0156 : integer;
		variable a0157 : integer;
		variable a0158 : integer;
		variable a0159 : integer;
		variable a0160 : integer;
		variable a0161 : integer;
		variable a0162 : integer;
		variable a0163 : integer;
		variable a0164 : integer;
		variable a0165 : integer;
		variable a0166 : integer;
		variable a0167 : integer;
		variable a0168 : integer;
		variable a0169 : integer;
		variable a0170 : integer;
		variable a0171 : integer;
		variable a0172 : integer;
		variable a0173 : integer;
		variable a0174 : integer;
		variable a0175 : integer;
		variable a0176 : integer;
		variable a0177 : integer;
		variable a0178 : integer;
		variable a0179 : integer;
		variable a0180 : integer;
		variable a0181 : integer;
		variable a0182 : integer;
		variable a0183 : integer;
		variable a0184 : integer;
		variable a0185 : integer;
		variable a0186 : integer;
		variable a0187 : integer;
		variable a0188 : integer;
		variable a0189 : integer;
		variable a0190 : integer;
		variable a0191 : integer;
		variable a0192 : integer;
		variable a0193 : integer;
		variable a0194 : integer;
		variable a0195 : integer;
		variable a0196 : integer;
		variable a0197 : integer;
		variable a0198 : integer;
		variable a0199 : integer;
		variable a0200 : integer;
		variable a0201 : integer;
		variable a0202 : integer;
		variable a0203 : integer;
		variable a0204 : integer;
		variable a0205 : integer;
		variable a0206 : integer;
		variable a0207 : integer;
		variable a0208 : integer;
		variable a0209 : integer;
		variable a0210 : integer;
		variable a0211 : integer;
		variable a0212 : integer;
		variable a0213 : integer;
		variable a0214 : integer;
		variable a0215 : integer;
		variable a0216 : integer;
		variable a0217 : integer;
		variable a0218 : integer;
		variable a0219 : integer;
		variable a0220 : integer;
		variable a0221 : integer;
		variable a0222 : integer;
		variable a0223 : integer;
		variable a0224 : integer;
		variable a0225 : integer;
		variable a0226 : integer;
		variable a0227 : integer;
		variable a0228 : integer;
		variable a0229 : integer;
		variable a0230 : integer;
		variable a0231 : integer;
		variable a0232 : integer;
		variable a0233 : integer;
		variable a0234 : integer;
		variable a0235 : integer;
		variable a0236 : integer;
		variable a0237 : integer;
		variable a0238 : integer;
		variable a0239 : integer;
		variable a0240 : integer;
		variable a0241 : integer;
		variable a0242 : integer;
		variable a0243 : integer;
		variable a0244 : integer;
		variable a0245 : integer;
		variable a0246 : integer;
		variable a0247 : integer;
		variable a0248 : integer;
		variable a0249 : integer;
		variable a0250 : integer;
		variable a0251 : integer;
		variable a0252 : integer;
		variable a0253 : integer;
		variable a0254 : integer;
		variable a0255 : integer;
		variable a0256 : integer;
		variable a0257 : integer;
		variable a0258 : integer;
		variable a0259 : integer;
		variable a0260 : integer;
		variable a0261 : integer;
		variable a0262 : integer;
		variable a0263 : integer;
		variable a0264 : integer;
		variable a0265 : integer;
		variable a0266 : integer;
		variable a0267 : integer;
		variable a0268 : integer;
		variable a0269 : integer;
		variable a0270 : integer;
		variable a0271 : integer;
		variable a0272 : integer;
		variable a0273 : integer;
		variable a0274 : integer;
		variable a0275 : integer;
		variable a0276 : integer;
		variable a0277 : integer;
		variable a0278 : integer;
		variable a0279 : integer;
		variable a0280 : integer;
		variable a0281 : integer;
		variable a0282 : integer;
		variable a0283 : integer;
		variable a0284 : integer;
		variable a0285 : integer;
		variable a0286 : integer;
		variable a0287 : integer;
		variable a0288 : integer;
		variable a0289 : integer;
		variable a0290 : integer;
		variable a0291 : integer;
		variable a0292 : integer;
		variable a0293 : integer;
		variable a0294 : integer;
		variable a0295 : integer;
		variable a0296 : integer;
		variable a0297 : integer;
		variable a0298 : integer;
		variable a0299 : integer;
		variable a0300 : integer;
		variable a0301 : integer;
		variable a0302 : integer;
		variable a0303 : integer;
		variable a0304 : integer;
		variable a0305 : integer;
		variable a0306 : integer;
		variable a0307 : integer;
		variable a0308 : integer;
		variable a0309 : integer;
		variable a0310 : integer;
		variable a0311 : integer;
		variable a0312 : integer;
		variable a0313 : integer;
		variable a0314 : integer;
		variable a0315 : integer;
		variable a0316 : integer;
		variable a0317 : integer;
		variable a0318 : integer;
		variable a0319 : integer;
		variable a0320 : integer;
		variable a0321 : integer;
		variable a0322 : integer;
		variable a0323 : integer;
		variable a0324 : integer;
		variable a0325 : integer;
		variable a0326 : integer;
		variable a0327 : integer;
		variable a0328 : integer;
		variable a0329 : integer;
		variable a0330 : integer;
		variable a0331 : integer;
		variable a0332 : integer;
		variable a0333 : integer;
		variable a0334 : integer;
		variable a0335 : integer;
		variable a0336 : integer;
		variable a0337 : integer;
		variable a0338 : integer;
		variable a0339 : integer;
		variable a0340 : integer;
		variable a0341 : integer;
		variable a0342 : integer;
		variable a0343 : integer;
		variable a0344 : integer;
		variable a0345 : integer;
		variable a0346 : integer;
		variable a0347 : integer;
		variable a0348 : integer;
		variable a0349 : integer;
		variable a0350 : integer;
		variable a0351 : integer;
		variable a0352 : integer;
		variable a0353 : integer;
		variable a0354 : integer;
		variable a0355 : integer;
		variable a0356 : integer;
		variable a0357 : integer;
		variable a0358 : integer;
		variable a0359 : integer;
		variable a0360 : integer;
		variable a0361 : integer;
		variable a0362 : integer;
		variable a0363 : integer;
		variable a0364 : integer;
		variable a0365 : integer;
		variable a0366 : integer;
		variable a0367 : integer;
		variable a0368 : integer;
		variable a0369 : integer;
		variable a0370 : integer;
		variable a0371 : integer;
		variable a0372 : integer;
		variable a0373 : integer;
		variable a0374 : integer;
		variable a0375 : integer;
		variable a0376 : integer;
		variable a0377 : integer;
		variable a0378 : integer;
		variable a0379 : integer;
		variable a0380 : integer;
		variable a0381 : integer;
		variable a0382 : integer;
		variable a0383 : integer;
		variable a0384 : integer;
		variable a0385 : integer;
		variable a0386 : integer;
		variable a0387 : integer;
		variable a0388 : integer;
		variable a0389 : integer;
		variable a0390 : integer;
		variable a0391 : integer;
		variable a0392 : integer;
		variable a0393 : integer;
		variable a0394 : integer;
		variable a0395 : integer;
		variable a0396 : integer;
		variable a0397 : integer;
		variable a0398 : integer;
		variable a0399 : integer;
		variable a0400 : integer;
		variable a0401 : integer;
		variable a0402 : integer;
		variable a0403 : integer;
		variable a0404 : integer;
		variable a0405 : integer;
		variable a0406 : integer;
		variable a0407 : integer;
		variable a0408 : integer;
		variable a0409 : integer;
		variable a0410 : integer;
		variable a0411 : integer;
		variable a0412 : integer;
		variable a0413 : integer;
		variable a0414 : integer;
		variable a0415 : integer;
		variable a0416 : integer;
		variable a0417 : integer;
		variable a0418 : integer;
		variable a0419 : integer;
		variable a0420 : integer;
		variable a0421 : integer;
		variable a0422 : integer;
		variable a0423 : integer;
		variable a0424 : integer;
		variable a0425 : integer;
		variable a0426 : integer;
		variable a0427 : integer;
		variable a0428 : integer;
		variable a0429 : integer;
		variable a0430 : integer;
		variable a0431 : integer;
		variable a0432 : integer;
		variable a0433 : integer;
		variable a0434 : integer;
		variable a0435 : integer;
		variable a0436 : integer;
		variable a0437 : integer;
		variable a0438 : integer;
		variable a0439 : integer;
		variable a0440 : integer;
		variable a0441 : integer;
		variable a0442 : integer;
		variable a0443 : integer;
		variable a0444 : integer;
		variable a0445 : integer;
		variable a0446 : integer;
		variable a0447 : integer;
		variable a0448 : integer;
		variable a0449 : integer;
		variable a0450 : integer;
		variable a0451 : integer;
		variable a0452 : integer;
		variable a0453 : integer;
		variable a0454 : integer;
		variable a0455 : integer;
		variable a0456 : integer;
		variable a0457 : integer;
		variable a0458 : integer;
		variable a0459 : integer;
		variable a0460 : integer;
		variable a0461 : integer;
		variable a0462 : integer;
		variable a0463 : integer;
		variable a0464 : integer;
		variable a0465 : integer;
		variable a0466 : integer;
		variable a0467 : integer;
		variable a0468 : integer;
		variable a0469 : integer;
		variable a0470 : integer;
		variable a0471 : integer;
		variable a0472 : integer;
		variable a0473 : integer;
		variable a0474 : integer;
		variable a0475 : integer;
		variable a0476 : integer;
		variable a0477 : integer;
		variable a0478 : integer;
		variable a0479 : integer;
		variable a0480 : integer;
		variable a0481 : integer;
		variable a0482 : integer;
		variable a0483 : integer;
		variable a0484 : integer;
		variable a0485 : integer;
		variable a0486 : integer;
		variable a0487 : integer;
		variable a0488 : integer;
		variable a0489 : integer;
		variable a0490 : integer;
		variable a0491 : integer;
		variable a0492 : integer;
		variable a0493 : integer;
		variable a0494 : integer;
		variable a0495 : integer;
		variable a0496 : integer;
		variable a0497 : integer;
		variable a0498 : integer;
		variable a0499 : integer;
		variable a0500 : integer;
		variable a0501 : integer;
		variable a0502 : integer;
		variable a0503 : integer;
		variable a0504 : integer;
		variable a0505 : integer;
		variable a0506 : integer;
		variable a0507 : integer;
		variable a0508 : integer;
		variable a0509 : integer;
		variable a0510 : integer;
		variable a0511 : integer;
		variable a0512 : integer;
		variable a0513 : integer;
		variable a0514 : integer;
		variable a0515 : integer;
		variable a0516 : integer;
		variable a0517 : integer;
		variable a0518 : integer;
		variable a0519 : integer;
		variable a0520 : integer;
		variable a0521 : integer;
		variable a0522 : integer;
		variable a0523 : integer;
		variable a0524 : integer;
		variable a0525 : integer;
		variable a0526 : integer;
		variable a0527 : integer;
		variable a0528 : integer;
		variable a0529 : integer;
		variable a0530 : integer;
		variable a0531 : integer;
		variable a0532 : integer;
		variable a0533 : integer;
		variable a0534 : integer;
		variable a0535 : integer;
		variable a0536 : integer;
		variable a0537 : integer;
		variable a0538 : integer;
		variable a0539 : integer;
		variable a0540 : integer;
		variable a0541 : integer;
		variable a0542 : integer;
		variable a0543 : integer;
		variable a0544 : integer;
		variable a0545 : integer;
		variable a0546 : integer;
		variable a0547 : integer;
		variable a0548 : integer;
		variable a0549 : integer;
		variable a0550 : integer;
		variable a0551 : integer;
		variable a0552 : integer;
		variable a0553 : integer;
		variable a0554 : integer;
		variable a0555 : integer;
		variable a0556 : integer;
		variable a0557 : integer;
		variable a0558 : integer;
		variable a0559 : integer;
		variable a0560 : integer;
		variable a0561 : integer;
		variable a0562 : integer;
		variable a0563 : integer;
		variable a0564 : integer;
		variable a0565 : integer;
		variable a0566 : integer;
		variable a0567 : integer;
		variable a0568 : integer;
		variable a0569 : integer;
		variable a0570 : integer;
		variable a0571 : integer;
		variable a0572 : integer;
		variable a0573 : integer;
		variable a0574 : integer;
		variable a0575 : integer;
		variable a0576 : integer;
		variable a0577 : integer;
		variable a0578 : integer;
		variable a0579 : integer;
		variable a0580 : integer;
		variable a0581 : integer;
		variable a0582 : integer;
		variable a0583 : integer;
		variable a0584 : integer;
		variable a0585 : integer;
		variable a0586 : integer;
		variable a0587 : integer;
		variable a0588 : integer;
		variable a0589 : integer;
		variable a0590 : integer;
		variable a0591 : integer;
		variable a0592 : integer;
		variable a0593 : integer;
		variable a0594 : integer;
		variable a0595 : integer;
		variable a0596 : integer;
		variable a0597 : integer;
		variable a0598 : integer;
		variable a0599 : integer;
		variable a0600 : integer;
		variable a0601 : integer;
		variable a0602 : integer;
		variable a0603 : integer;
		variable a0604 : integer;
		variable a0605 : integer;
		variable a0606 : integer;
		variable a0607 : integer;
		variable a0608 : integer;
		variable a0609 : integer;
		variable a0610 : integer;
		variable a0611 : integer;
		variable a0612 : integer;
		variable a0613 : integer;
		variable a0614 : integer;
		variable a0615 : integer;
		variable a0616 : integer;
		variable a0617 : integer;
		variable a0618 : integer;
		variable a0619 : integer;
		variable a0620 : integer;
		variable a0621 : integer;
		variable a0622 : integer;
		variable a0623 : integer;
		variable a0624 : integer;
		variable a0625 : integer;
		variable a0626 : integer;
		variable a0627 : integer;
		variable a0628 : integer;
		variable a0629 : integer;
		variable a0630 : integer;
		variable a0631 : integer;
		variable a0632 : integer;
		variable a0633 : integer;
		variable a0634 : integer;
		variable a0635 : integer;
		variable a0636 : integer;
		variable a0637 : integer;
		variable a0638 : integer;
		variable a0639 : integer;
		variable a0640 : integer;
		variable a0641 : integer;
		variable a0642 : integer;
		variable a0643 : integer;
		variable a0644 : integer;
		variable a0645 : integer;
		variable a0646 : integer;
		variable a0647 : integer;
		variable a0648 : integer;
		variable a0649 : integer;
		variable a0650 : integer;
		variable a0651 : integer;
		variable a0652 : integer;
		variable a0653 : integer;
		variable a0654 : integer;
		variable a0655 : integer;
		variable a0656 : integer;
		variable a0657 : integer;
		variable a0658 : integer;
		variable a0659 : integer;
		variable a0660 : integer;
		variable a0661 : integer;
		variable a0662 : integer;
		variable a0663 : integer;
		variable a0664 : integer;
		variable a0665 : integer;
		variable a0666 : integer;
		variable a0667 : integer;
		variable a0668 : integer;
		variable a0669 : integer;
		variable a0670 : integer;
		variable a0671 : integer;
		variable a0672 : integer;
		variable a0673 : integer;
		variable a0674 : integer;
		variable a0675 : integer;
		variable a0676 : integer;
		variable a0677 : integer;
		variable a0678 : integer;
		variable a0679 : integer;
		variable a0680 : integer;
		variable a0681 : integer;
		variable a0682 : integer;
		variable a0683 : integer;
		variable a0684 : integer;
		variable a0685 : integer;
		variable a0686 : integer;
		variable a0687 : integer;
		variable a0688 : integer;
		variable a0689 : integer;
		variable a0690 : integer;
		variable a0691 : integer;
		variable a0692 : integer;
		variable a0693 : integer;
		variable a0694 : integer;
		variable a0695 : integer;
		variable a0696 : integer;
		variable a0697 : integer;
		variable a0698 : integer;
		variable a0699 : integer;
		variable a0700 : integer;
		variable a0701 : integer;
		variable a0702 : integer;
		variable a0703 : integer;
		variable a0704 : integer;
		variable a0705 : integer;
		variable a0706 : integer;
		variable a0707 : integer;
		variable a0708 : integer;
		variable a0709 : integer;
		variable a0710 : integer;
		variable a0711 : integer;
		variable a0712 : integer;
		variable a0713 : integer;
		variable a0714 : integer;
		variable a0715 : integer;
		variable a0716 : integer;
		variable a0717 : integer;
		variable a0718 : integer;
		variable a0719 : integer;
		variable a0720 : integer;
		variable a0721 : integer;
		variable a0722 : integer;
		variable a0723 : integer;
		variable a0724 : integer;
		variable a0725 : integer;
		variable a0726 : integer;
		variable a0727 : integer;
		variable a0728 : integer;
		variable a0729 : integer;
		variable a0730 : integer;
		variable a0731 : integer;
		variable a0732 : integer;
		variable a0733 : integer;
		variable a0734 : integer;
		variable a0735 : integer;
		variable a0736 : integer;
		variable a0737 : integer;
		variable a0738 : integer;
		variable a0739 : integer;
		variable a0740 : integer;
		variable a0741 : integer;
		variable a0742 : integer;
		variable a0743 : integer;
		variable a0744 : integer;
		variable a0745 : integer;
		variable a0746 : integer;
		variable a0747 : integer;
		variable a0748 : integer;
		variable a0749 : integer;
		variable a0750 : integer;
		variable a0751 : integer;
		variable a0752 : integer;
		variable a0753 : integer;
		variable a0754 : integer;
		variable a0755 : integer;
		variable a0756 : integer;
		variable a0757 : integer;
		variable a0758 : integer;
		variable a0759 : integer;
		variable a0760 : integer;
		variable a0761 : integer;
		variable a0762 : integer;
		variable a0763 : integer;
		variable a0764 : integer;
		variable a0765 : integer;
		variable a0766 : integer;
		variable a0767 : integer;
		variable a0768 : integer;
		variable a0769 : integer;
		variable a0770 : integer;
		variable a0771 : integer;
		variable a0772 : integer;
		variable a0773 : integer;
		variable a0774 : integer;
		variable a0775 : integer;
		variable a0776 : integer;
		variable a0777 : integer;
		variable a0778 : integer;
		variable a0779 : integer;
		variable a0780 : integer;
		variable a0781 : integer;
		variable a0782 : integer;
		variable a0783 : integer;
		variable a0784 : integer;
		variable a0785 : integer;
		variable a0786 : integer;
		variable a0787 : integer;
		variable a0788 : integer;
		variable a0789 : integer;
		variable a0790 : integer;
		variable a0791 : integer;
		variable a0792 : integer;
		variable a0793 : integer;
		variable a0794 : integer;
		variable a0795 : integer;
		variable a0796 : integer;
		variable a0797 : integer;
		variable a0798 : integer;
		variable a0799 : integer;
		variable a0800 : integer;
		variable a0801 : integer;
		variable a0802 : integer;
		variable a0803 : integer;
		variable a0804 : integer;
		variable a0805 : integer;
		variable a0806 : integer;
		variable a0807 : integer;
		variable a0808 : integer;
		variable a0809 : integer;
		variable a0810 : integer;
		variable a0811 : integer;
		variable a0812 : integer;
		variable a0813 : integer;
		variable a0814 : integer;
		variable a0815 : integer;
		variable a0816 : integer;
		variable a0817 : integer;
		variable a0818 : integer;
		variable a0819 : integer;
		variable a0820 : integer;
		variable a0821 : integer;
		variable a0822 : integer;
		variable a0823 : integer;
		variable a0824 : integer;
		variable a0825 : integer;
		variable a0826 : integer;
		variable a0827 : integer;
		variable a0828 : integer;
		variable a0829 : integer;
		variable a0830 : integer;
		variable a0831 : integer;
		variable a0832 : integer;
		variable a0833 : integer;
		variable a0834 : integer;
		variable a0835 : integer;
		variable a0836 : integer;
		variable a0837 : integer;
		variable a0838 : integer;
		variable a0839 : integer;
		variable a0840 : integer;
		variable a0841 : integer;
		variable a0842 : integer;
		variable a0843 : integer;
		variable a0844 : integer;
		variable a0845 : integer;
		variable a0846 : integer;
		variable a0847 : integer;
		variable a0848 : integer;
		variable a0849 : integer;
		variable a0850 : integer;
		variable a0851 : integer;
		variable a0852 : integer;
		variable a0853 : integer;
		variable a0854 : integer;
		variable a0855 : integer;
		variable a0856 : integer;
		variable a0857 : integer;
		variable a0858 : integer;
		variable a0859 : integer;
		variable a0860 : integer;
		variable a0861 : integer;
		variable a0862 : integer;
		variable a0863 : integer;
		variable a0864 : integer;
		variable a0865 : integer;
		variable a0866 : integer;
		variable a0867 : integer;
		variable a0868 : integer;
		variable a0869 : integer;
		variable a0870 : integer;
		variable a0871 : integer;
		variable a0872 : integer;
		variable a0873 : integer;
		variable a0874 : integer;
		variable a0875 : integer;
		variable a0876 : integer;
		variable a0877 : integer;
		variable a0878 : integer;
		variable a0879 : integer;
		variable a0880 : integer;
		variable a0881 : integer;
		variable a0882 : integer;
		variable a0883 : integer;
		variable a0884 : integer;
		variable a0885 : integer;
		variable a0886 : integer;
		variable a0887 : integer;
		variable a0888 : integer;
		variable a0889 : integer;
		variable a0890 : integer;
		variable a0891 : integer;
		variable a0892 : integer;
		variable a0893 : integer;
		variable a0894 : integer;
		variable a0895 : integer;
		variable a0896 : integer;
		variable a0897 : integer;
		variable a0898 : integer;
		variable a0899 : integer;
		variable a0900 : integer;
		variable a0901 : integer;
		variable a0902 : integer;
		variable a0903 : integer;
		variable a0904 : integer;
		variable a0905 : integer;
		variable a0906 : integer;
		variable a0907 : integer;
		variable a0908 : integer;
		variable a0909 : integer;
		variable a0910 : integer;
		variable a0911 : integer;
		variable a0912 : integer;
		variable a0913 : integer;
		variable a0914 : integer;
		variable a0915 : integer;
		variable a0916 : integer;
		variable a0917 : integer;
		variable a0918 : integer;
		variable a0919 : integer;
		variable a0920 : integer;
		variable a0921 : integer;
		variable a0922 : integer;
		variable a0923 : integer;
		variable a0924 : integer;
		variable a0925 : integer;
		variable a0926 : integer;
		variable a0927 : integer;
		variable a0928 : integer;
		variable a0929 : integer;
		variable a0930 : integer;
		variable a0931 : integer;
		variable a0932 : integer;
		variable a0933 : integer;
		variable a0934 : integer;
		variable a0935 : integer;
		variable a0936 : integer;
		variable a0937 : integer;
		variable a0938 : integer;
		variable a0939 : integer;
		variable a0940 : integer;
		variable a0941 : integer;
		variable a0942 : integer;
		variable a0943 : integer;
		variable a0944 : integer;
		variable a0945 : integer;
		variable a0946 : integer;
		variable a0947 : integer;
		variable a0948 : integer;
		variable a0949 : integer;
		variable a0950 : integer;
		variable a0951 : integer;
		variable a0952 : integer;
		variable a0953 : integer;
		variable a0954 : integer;
		variable a0955 : integer;
		variable a0956 : integer;
		variable a0957 : integer;
		variable a0958 : integer;
		variable a0959 : integer;
		variable a0960 : integer;
		variable a0961 : integer;
		variable a0962 : integer;
		variable a0963 : integer;
		variable a0964 : integer;
		variable a0965 : integer;
		variable a0966 : integer;
		variable a0967 : integer;
		variable a0968 : integer;
		variable a0969 : integer;
		variable a0970 : integer;
		variable a0971 : integer;
		variable a0972 : integer;
		variable a0973 : integer;
		variable a0974 : integer;
		variable a0975 : integer;
		variable a0976 : integer;
		variable a0977 : integer;
		variable a0978 : integer;
		variable a0979 : integer;
		variable a0980 : integer;
		variable a0981 : integer;
		variable a0982 : integer;
		variable a0983 : integer;
		variable a0984 : integer;
		variable a0985 : integer;
		variable a0986 : integer;
		variable a0987 : integer;
		variable a0988 : integer;
		variable a0989 : integer;
		variable a0990 : integer;
		variable a0991 : integer;
		variable a0992 : integer;
		variable a0993 : integer;
		variable a0994 : integer;
		variable a0995 : integer;
		variable a0996 : integer;
		variable a0997 : integer;
		variable a0998 : integer;
		variable a0999 : integer;
		variable a1000 : integer;
	begin

		a0001 := clk;
		a0002 := clk;
		a0003 := clk;
		a0004 := clk;
		a0005 := clk;
		a0006 := clk;
		a0007 := clk;
		a0008 := clk;
		a0009 := clk;
		a0010 := clk;
		a0011 := clk;
		a0012 := clk;
		a0013 := clk;
		a0014 := clk;
		a0015 := clk;
		a0016 := clk;
		a0017 := clk;
		a0018 := clk;
		a0019 := clk;
		a0020 := clk;
		a0021 := clk;
		a0022 := clk;
		a0023 := clk;
		a0024 := clk;
		a0025 := clk;
		a0026 := clk;
		a0027 := clk;
		a0028 := clk;
		a0029 := clk;
		a0030 := clk;
		a0031 := clk;
		a0032 := clk;
		a0033 := clk;
		a0034 := clk;
		a0035 := clk;
		a0036 := clk;
		a0037 := clk;
		a0038 := clk;
		a0039 := clk;
		a0040 := clk;
		a0041 := clk;
		a0042 := clk;
		a0043 := clk;
		a0044 := clk;
		a0045 := clk;
		a0046 := clk;
		a0047 := clk;
		a0048 := clk;
		a0049 := clk;
		a0050 := clk;
		a0051 := clk;
		a0052 := clk;
		a0053 := clk;
		a0054 := clk;
		a0055 := clk;
		a0056 := clk;
		a0057 := clk;
		a0058 := clk;
		a0059 := clk;
		a0060 := clk;
		a0061 := clk;
		a0062 := clk;
		a0063 := clk;
		a0064 := clk;
		a0065 := clk;
		a0066 := clk;
		a0067 := clk;
		a0068 := clk;
		a0069 := clk;
		a0070 := clk;
		a0071 := clk;
		a0072 := clk;
		a0073 := clk;
		a0074 := clk;
		a0075 := clk;
		a0076 := clk;
		a0077 := clk;
		a0078 := clk;
		a0079 := clk;
		a0080 := clk;
		a0081 := clk;
		a0082 := clk;
		a0083 := clk;
		a0084 := clk;
		a0085 := clk;
		a0086 := clk;
		a0087 := clk;
		a0088 := clk;
		a0089 := clk;
		a0090 := clk;
		a0091 := clk;
		a0092 := clk;
		a0093 := clk;
		a0094 := clk;
		a0095 := clk;
		a0096 := clk;
		a0097 := clk;
		a0098 := clk;
		a0099 := clk;
		a0100 := clk;
		a0101 := clk;
		a0102 := clk;
		a0103 := clk;
		a0104 := clk;
		a0105 := clk;
		a0106 := clk;
		a0107 := clk;
		a0108 := clk;
		a0109 := clk;
		a0110 := clk;
		a0111 := clk;
		a0112 := clk;
		a0113 := clk;
		a0114 := clk;
		a0115 := clk;
		a0116 := clk;
		a0117 := clk;
		a0118 := clk;
		a0119 := clk;
		a0120 := clk;
		a0121 := clk;
		a0122 := clk;
		a0123 := clk;
		a0124 := clk;
		a0125 := clk;
		a0126 := clk;
		a0127 := clk;
		a0128 := clk;
		a0129 := clk;
		a0130 := clk;
		a0131 := clk;
		a0132 := clk;
		a0133 := clk;
		a0134 := clk;
		a0135 := clk;
		a0136 := clk;
		a0137 := clk;
		a0138 := clk;
		a0139 := clk;
		a0140 := clk;
		a0141 := clk;
		a0142 := clk;
		a0143 := clk;
		a0144 := clk;
		a0145 := clk;
		a0146 := clk;
		a0147 := clk;
		a0148 := clk;
		a0149 := clk;
		a0150 := clk;
		a0151 := clk;
		a0152 := clk;
		a0153 := clk;
		a0154 := clk;
		a0155 := clk;
		a0156 := clk;
		a0157 := clk;
		a0158 := clk;
		a0159 := clk;
		a0160 := clk;
		a0161 := clk;
		a0162 := clk;
		a0163 := clk;
		a0164 := clk;
		a0165 := clk;
		a0166 := clk;
		a0167 := clk;
		a0168 := clk;
		a0169 := clk;
		a0170 := clk;
		a0171 := clk;
		a0172 := clk;
		a0173 := clk;
		a0174 := clk;
		a0175 := clk;
		a0176 := clk;
		a0177 := clk;
		a0178 := clk;
		a0179 := clk;
		a0180 := clk;
		a0181 := clk;
		a0182 := clk;
		a0183 := clk;
		a0184 := clk;
		a0185 := clk;
		a0186 := clk;
		a0187 := clk;
		a0188 := clk;
		a0189 := clk;
		a0190 := clk;
		a0191 := clk;
		a0192 := clk;
		a0193 := clk;
		a0194 := clk;
		a0195 := clk;
		a0196 := clk;
		a0197 := clk;
		a0198 := clk;
		a0199 := clk;
		a0200 := clk;
		a0201 := clk;
		a0202 := clk;
		a0203 := clk;
		a0204 := clk;
		a0205 := clk;
		a0206 := clk;
		a0207 := clk;
		a0208 := clk;
		a0209 := clk;
		a0210 := clk;
		a0211 := clk;
		a0212 := clk;
		a0213 := clk;
		a0214 := clk;
		a0215 := clk;
		a0216 := clk;
		a0217 := clk;
		a0218 := clk;
		a0219 := clk;
		a0220 := clk;
		a0221 := clk;
		a0222 := clk;
		a0223 := clk;
		a0224 := clk;
		a0225 := clk;
		a0226 := clk;
		a0227 := clk;
		a0228 := clk;
		a0229 := clk;
		a0230 := clk;
		a0231 := clk;
		a0232 := clk;
		a0233 := clk;
		a0234 := clk;
		a0235 := clk;
		a0236 := clk;
		a0237 := clk;
		a0238 := clk;
		a0239 := clk;
		a0240 := clk;
		a0241 := clk;
		a0242 := clk;
		a0243 := clk;
		a0244 := clk;
		a0245 := clk;
		a0246 := clk;
		a0247 := clk;
		a0248 := clk;
		a0249 := clk;
		a0250 := clk;
		a0251 := clk;
		a0252 := clk;
		a0253 := clk;
		a0254 := clk;
		a0255 := clk;
		a0256 := clk;
		a0257 := clk;
		a0258 := clk;
		a0259 := clk;
		a0260 := clk;
		a0261 := clk;
		a0262 := clk;
		a0263 := clk;
		a0264 := clk;
		a0265 := clk;
		a0266 := clk;
		a0267 := clk;
		a0268 := clk;
		a0269 := clk;
		a0270 := clk;
		a0271 := clk;
		a0272 := clk;
		a0273 := clk;
		a0274 := clk;
		a0275 := clk;
		a0276 := clk;
		a0277 := clk;
		a0278 := clk;
		a0279 := clk;
		a0280 := clk;
		a0281 := clk;
		a0282 := clk;
		a0283 := clk;
		a0284 := clk;
		a0285 := clk;
		a0286 := clk;
		a0287 := clk;
		a0288 := clk;
		a0289 := clk;
		a0290 := clk;
		a0291 := clk;
		a0292 := clk;
		a0293 := clk;
		a0294 := clk;
		a0295 := clk;
		a0296 := clk;
		a0297 := clk;
		a0298 := clk;
		a0299 := clk;
		a0300 := clk;
		a0301 := clk;
		a0302 := clk;
		a0303 := clk;
		a0304 := clk;
		a0305 := clk;
		a0306 := clk;
		a0307 := clk;
		a0308 := clk;
		a0309 := clk;
		a0310 := clk;
		a0311 := clk;
		a0312 := clk;
		a0313 := clk;
		a0314 := clk;
		a0315 := clk;
		a0316 := clk;
		a0317 := clk;
		a0318 := clk;
		a0319 := clk;
		a0320 := clk;
		a0321 := clk;
		a0322 := clk;
		a0323 := clk;
		a0324 := clk;
		a0325 := clk;
		a0326 := clk;
		a0327 := clk;
		a0328 := clk;
		a0329 := clk;
		a0330 := clk;
		a0331 := clk;
		a0332 := clk;
		a0333 := clk;
		a0334 := clk;
		a0335 := clk;
		a0336 := clk;
		a0337 := clk;
		a0338 := clk;
		a0339 := clk;
		a0340 := clk;
		a0341 := clk;
		a0342 := clk;
		a0343 := clk;
		a0344 := clk;
		a0345 := clk;
		a0346 := clk;
		a0347 := clk;
		a0348 := clk;
		a0349 := clk;
		a0350 := clk;
		a0351 := clk;
		a0352 := clk;
		a0353 := clk;
		a0354 := clk;
		a0355 := clk;
		a0356 := clk;
		a0357 := clk;
		a0358 := clk;
		a0359 := clk;
		a0360 := clk;
		a0361 := clk;
		a0362 := clk;
		a0363 := clk;
		a0364 := clk;
		a0365 := clk;
		a0366 := clk;
		a0367 := clk;
		a0368 := clk;
		a0369 := clk;
		a0370 := clk;
		a0371 := clk;
		a0372 := clk;
		a0373 := clk;
		a0374 := clk;
		a0375 := clk;
		a0376 := clk;
		a0377 := clk;
		a0378 := clk;
		a0379 := clk;
		a0380 := clk;
		a0381 := clk;
		a0382 := clk;
		a0383 := clk;
		a0384 := clk;
		a0385 := clk;
		a0386 := clk;
		a0387 := clk;
		a0388 := clk;
		a0389 := clk;
		a0390 := clk;
		a0391 := clk;
		a0392 := clk;
		a0393 := clk;
		a0394 := clk;
		a0395 := clk;
		a0396 := clk;
		a0397 := clk;
		a0398 := clk;
		a0399 := clk;
		a0400 := clk;
		a0401 := clk;
		a0402 := clk;
		a0403 := clk;
		a0404 := clk;
		a0405 := clk;
		a0406 := clk;
		a0407 := clk;
		a0408 := clk;
		a0409 := clk;
		a0410 := clk;
		a0411 := clk;
		a0412 := clk;
		a0413 := clk;
		a0414 := clk;
		a0415 := clk;
		a0416 := clk;
		a0417 := clk;
		a0418 := clk;
		a0419 := clk;
		a0420 := clk;
		a0421 := clk;
		a0422 := clk;
		a0423 := clk;
		a0424 := clk;
		a0425 := clk;
		a0426 := clk;
		a0427 := clk;
		a0428 := clk;
		a0429 := clk;
		a0430 := clk;
		a0431 := clk;
		a0432 := clk;
		a0433 := clk;
		a0434 := clk;
		a0435 := clk;
		a0436 := clk;
		a0437 := clk;
		a0438 := clk;
		a0439 := clk;
		a0440 := clk;
		a0441 := clk;
		a0442 := clk;
		a0443 := clk;
		a0444 := clk;
		a0445 := clk;
		a0446 := clk;
		a0447 := clk;
		a0448 := clk;
		a0449 := clk;
		a0450 := clk;
		a0451 := clk;
		a0452 := clk;
		a0453 := clk;
		a0454 := clk;
		a0455 := clk;
		a0456 := clk;
		a0457 := clk;
		a0458 := clk;
		a0459 := clk;
		a0460 := clk;
		a0461 := clk;
		a0462 := clk;
		a0463 := clk;
		a0464 := clk;
		a0465 := clk;
		a0466 := clk;
		a0467 := clk;
		a0468 := clk;
		a0469 := clk;
		a0470 := clk;
		a0471 := clk;
		a0472 := clk;
		a0473 := clk;
		a0474 := clk;
		a0475 := clk;
		a0476 := clk;
		a0477 := clk;
		a0478 := clk;
		a0479 := clk;
		a0480 := clk;
		a0481 := clk;
		a0482 := clk;
		a0483 := clk;
		a0484 := clk;
		a0485 := clk;
		a0486 := clk;
		a0487 := clk;
		a0488 := clk;
		a0489 := clk;
		a0490 := clk;
		a0491 := clk;
		a0492 := clk;
		a0493 := clk;
		a0494 := clk;
		a0495 := clk;
		a0496 := clk;
		a0497 := clk;
		a0498 := clk;
		a0499 := clk;
		a0500 := clk;
		a0501 := clk;
		a0502 := clk;
		a0503 := clk;
		a0504 := clk;
		a0505 := clk;
		a0506 := clk;
		a0507 := clk;
		a0508 := clk;
		a0509 := clk;
		a0510 := clk;
		a0511 := clk;
		a0512 := clk;
		a0513 := clk;
		a0514 := clk;
		a0515 := clk;
		a0516 := clk;
		a0517 := clk;
		a0518 := clk;
		a0519 := clk;
		a0520 := clk;
		a0521 := clk;
		a0522 := clk;
		a0523 := clk;
		a0524 := clk;
		a0525 := clk;
		a0526 := clk;
		a0527 := clk;
		a0528 := clk;
		a0529 := clk;
		a0530 := clk;
		a0531 := clk;
		a0532 := clk;
		a0533 := clk;
		a0534 := clk;
		a0535 := clk;
		a0536 := clk;
		a0537 := clk;
		a0538 := clk;
		a0539 := clk;
		a0540 := clk;
		a0541 := clk;
		a0542 := clk;
		a0543 := clk;
		a0544 := clk;
		a0545 := clk;
		a0546 := clk;
		a0547 := clk;
		a0548 := clk;
		a0549 := clk;
		a0550 := clk;
		a0551 := clk;
		a0552 := clk;
		a0553 := clk;
		a0554 := clk;
		a0555 := clk;
		a0556 := clk;
		a0557 := clk;
		a0558 := clk;
		a0559 := clk;
		a0560 := clk;
		a0561 := clk;
		a0562 := clk;
		a0563 := clk;
		a0564 := clk;
		a0565 := clk;
		a0566 := clk;
		a0567 := clk;
		a0568 := clk;
		a0569 := clk;
		a0570 := clk;
		a0571 := clk;
		a0572 := clk;
		a0573 := clk;
		a0574 := clk;
		a0575 := clk;
		a0576 := clk;
		a0577 := clk;
		a0578 := clk;
		a0579 := clk;
		a0580 := clk;
		a0581 := clk;
		a0582 := clk;
		a0583 := clk;
		a0584 := clk;
		a0585 := clk;
		a0586 := clk;
		a0587 := clk;
		a0588 := clk;
		a0589 := clk;
		a0590 := clk;
		a0591 := clk;
		a0592 := clk;
		a0593 := clk;
		a0594 := clk;
		a0595 := clk;
		a0596 := clk;
		a0597 := clk;
		a0598 := clk;
		a0599 := clk;
		a0600 := clk;
		a0601 := clk;
		a0602 := clk;
		a0603 := clk;
		a0604 := clk;
		a0605 := clk;
		a0606 := clk;
		a0607 := clk;
		a0608 := clk;
		a0609 := clk;
		a0610 := clk;
		a0611 := clk;
		a0612 := clk;
		a0613 := clk;
		a0614 := clk;
		a0615 := clk;
		a0616 := clk;
		a0617 := clk;
		a0618 := clk;
		a0619 := clk;
		a0620 := clk;
		a0621 := clk;
		a0622 := clk;
		a0623 := clk;
		a0624 := clk;
		a0625 := clk;
		a0626 := clk;
		a0627 := clk;
		a0628 := clk;
		a0629 := clk;
		a0630 := clk;
		a0631 := clk;
		a0632 := clk;
		a0633 := clk;
		a0634 := clk;
		a0635 := clk;
		a0636 := clk;
		a0637 := clk;
		a0638 := clk;
		a0639 := clk;
		a0640 := clk;
		a0641 := clk;
		a0642 := clk;
		a0643 := clk;
		a0644 := clk;
		a0645 := clk;
		a0646 := clk;
		a0647 := clk;
		a0648 := clk;
		a0649 := clk;
		a0650 := clk;
		a0651 := clk;
		a0652 := clk;
		a0653 := clk;
		a0654 := clk;
		a0655 := clk;
		a0656 := clk;
		a0657 := clk;
		a0658 := clk;
		a0659 := clk;
		a0660 := clk;
		a0661 := clk;
		a0662 := clk;
		a0663 := clk;
		a0664 := clk;
		a0665 := clk;
		a0666 := clk;
		a0667 := clk;
		a0668 := clk;
		a0669 := clk;
		a0670 := clk;
		a0671 := clk;
		a0672 := clk;
		a0673 := clk;
		a0674 := clk;
		a0675 := clk;
		a0676 := clk;
		a0677 := clk;
		a0678 := clk;
		a0679 := clk;
		a0680 := clk;
		a0681 := clk;
		a0682 := clk;
		a0683 := clk;
		a0684 := clk;
		a0685 := clk;
		a0686 := clk;
		a0687 := clk;
		a0688 := clk;
		a0689 := clk;
		a0690 := clk;
		a0691 := clk;
		a0692 := clk;
		a0693 := clk;
		a0694 := clk;
		a0695 := clk;
		a0696 := clk;
		a0697 := clk;
		a0698 := clk;
		a0699 := clk;
		a0700 := clk;
		a0701 := clk;
		a0702 := clk;
		a0703 := clk;
		a0704 := clk;
		a0705 := clk;
		a0706 := clk;
		a0707 := clk;
		a0708 := clk;
		a0709 := clk;
		a0710 := clk;
		a0711 := clk;
		a0712 := clk;
		a0713 := clk;
		a0714 := clk;
		a0715 := clk;
		a0716 := clk;
		a0717 := clk;
		a0718 := clk;
		a0719 := clk;
		a0720 := clk;
		a0721 := clk;
		a0722 := clk;
		a0723 := clk;
		a0724 := clk;
		a0725 := clk;
		a0726 := clk;
		a0727 := clk;
		a0728 := clk;
		a0729 := clk;
		a0730 := clk;
		a0731 := clk;
		a0732 := clk;
		a0733 := clk;
		a0734 := clk;
		a0735 := clk;
		a0736 := clk;
		a0737 := clk;
		a0738 := clk;
		a0739 := clk;
		a0740 := clk;
		a0741 := clk;
		a0742 := clk;
		a0743 := clk;
		a0744 := clk;
		a0745 := clk;
		a0746 := clk;
		a0747 := clk;
		a0748 := clk;
		a0749 := clk;
		a0750 := clk;
		a0751 := clk;
		a0752 := clk;
		a0753 := clk;
		a0754 := clk;
		a0755 := clk;
		a0756 := clk;
		a0757 := clk;
		a0758 := clk;
		a0759 := clk;
		a0760 := clk;
		a0761 := clk;
		a0762 := clk;
		a0763 := clk;
		a0764 := clk;
		a0765 := clk;
		a0766 := clk;
		a0767 := clk;
		a0768 := clk;
		a0769 := clk;
		a0770 := clk;
		a0771 := clk;
		a0772 := clk;
		a0773 := clk;
		a0774 := clk;
		a0775 := clk;
		a0776 := clk;
		a0777 := clk;
		a0778 := clk;
		a0779 := clk;
		a0780 := clk;
		a0781 := clk;
		a0782 := clk;
		a0783 := clk;
		a0784 := clk;
		a0785 := clk;
		a0786 := clk;
		a0787 := clk;
		a0788 := clk;
		a0789 := clk;
		a0790 := clk;
		a0791 := clk;
		a0792 := clk;
		a0793 := clk;
		a0794 := clk;
		a0795 := clk;
		a0796 := clk;
		a0797 := clk;
		a0798 := clk;
		a0799 := clk;
		a0800 := clk;
		a0801 := clk;
		a0802 := clk;
		a0803 := clk;
		a0804 := clk;
		a0805 := clk;
		a0806 := clk;
		a0807 := clk;
		a0808 := clk;
		a0809 := clk;
		a0810 := clk;
		a0811 := clk;
		a0812 := clk;
		a0813 := clk;
		a0814 := clk;
		a0815 := clk;
		a0816 := clk;
		a0817 := clk;
		a0818 := clk;
		a0819 := clk;
		a0820 := clk;
		a0821 := clk;
		a0822 := clk;
		a0823 := clk;
		a0824 := clk;
		a0825 := clk;
		a0826 := clk;
		a0827 := clk;
		a0828 := clk;
		a0829 := clk;
		a0830 := clk;
		a0831 := clk;
		a0832 := clk;
		a0833 := clk;
		a0834 := clk;
		a0835 := clk;
		a0836 := clk;
		a0837 := clk;
		a0838 := clk;
		a0839 := clk;
		a0840 := clk;
		a0841 := clk;
		a0842 := clk;
		a0843 := clk;
		a0844 := clk;
		a0845 := clk;
		a0846 := clk;
		a0847 := clk;
		a0848 := clk;
		a0849 := clk;
		a0850 := clk;
		a0851 := clk;
		a0852 := clk;
		a0853 := clk;
		a0854 := clk;
		a0855 := clk;
		a0856 := clk;
		a0857 := clk;
		a0858 := clk;
		a0859 := clk;
		a0860 := clk;
		a0861 := clk;
		a0862 := clk;
		a0863 := clk;
		a0864 := clk;
		a0865 := clk;
		a0866 := clk;
		a0867 := clk;
		a0868 := clk;
		a0869 := clk;
		a0870 := clk;
		a0871 := clk;
		a0872 := clk;
		a0873 := clk;
		a0874 := clk;
		a0875 := clk;
		a0876 := clk;
		a0877 := clk;
		a0878 := clk;
		a0879 := clk;
		a0880 := clk;
		a0881 := clk;
		a0882 := clk;
		a0883 := clk;
		a0884 := clk;
		a0885 := clk;
		a0886 := clk;
		a0887 := clk;
		a0888 := clk;
		a0889 := clk;
		a0890 := clk;
		a0891 := clk;
		a0892 := clk;
		a0893 := clk;
		a0894 := clk;
		a0895 := clk;
		a0896 := clk;
		a0897 := clk;
		a0898 := clk;
		a0899 := clk;
		a0900 := clk;
		a0901 := clk;
		a0902 := clk;
		a0903 := clk;
		a0904 := clk;
		a0905 := clk;
		a0906 := clk;
		a0907 := clk;
		a0908 := clk;
		a0909 := clk;
		a0910 := clk;
		a0911 := clk;
		a0912 := clk;
		a0913 := clk;
		a0914 := clk;
		a0915 := clk;
		a0916 := clk;
		a0917 := clk;
		a0918 := clk;
		a0919 := clk;
		a0920 := clk;
		a0921 := clk;
		a0922 := clk;
		a0923 := clk;
		a0924 := clk;
		a0925 := clk;
		a0926 := clk;
		a0927 := clk;
		a0928 := clk;
		a0929 := clk;
		a0930 := clk;
		a0931 := clk;
		a0932 := clk;
		a0933 := clk;
		a0934 := clk;
		a0935 := clk;
		a0936 := clk;
		a0937 := clk;
		a0938 := clk;
		a0939 := clk;
		a0940 := clk;
		a0941 := clk;
		a0942 := clk;
		a0943 := clk;
		a0944 := clk;
		a0945 := clk;
		a0946 := clk;
		a0947 := clk;
		a0948 := clk;
		a0949 := clk;
		a0950 := clk;
		a0951 := clk;
		a0952 := clk;
		a0953 := clk;
		a0954 := clk;
		a0955 := clk;
		a0956 := clk;
		a0957 := clk;
		a0958 := clk;
		a0959 := clk;
		a0960 := clk;
		a0961 := clk;
		a0962 := clk;
		a0963 := clk;
		a0964 := clk;
		a0965 := clk;
		a0966 := clk;
		a0967 := clk;
		a0968 := clk;
		a0969 := clk;
		a0970 := clk;
		a0971 := clk;
		a0972 := clk;
		a0973 := clk;
		a0974 := clk;
		a0975 := clk;
		a0976 := clk;
		a0977 := clk;
		a0978 := clk;
		a0979 := clk;
		a0980 := clk;
		a0981 := clk;
		a0982 := clk;
		a0983 := clk;
		a0984 := clk;
		a0985 := clk;
		a0986 := clk;
		a0987 := clk;
		a0988 := clk;
		a0989 := clk;
		a0990 := clk;
		a0991 := clk;
		a0992 := clk;
		a0993 := clk;
		a0994 := clk;
		a0995 := clk;
		a0996 := clk;
		a0997 := clk;
		a0998 := clk;
		a0999 := clk;
		a1000 := clk;
--}}}
    end process;

	terminator : process(clk)
	begin
		if clk >= CYCLES then
			assert false report "end of simulation" severity failure;
		-- else
		-- 	report "tick";
		end if;
	end process;

	clk <= (clk+1) after 1 us;
end;
