-- NEED RESULT: ENT00703: Open composite buffer ports with static subtypes passed
-------------------------------------------------------------------------------
 --
 --    Copyright (c) 1989 by Intermetrics, Inc.
 --                All rights reserved.
 --
-------------------------------------------------------------------------------
--
-- TEST NAME:
--
--    CT00703
--
-- AUTHOR:
--
--    A. Wilmot
--
-- TEST OBJECTIVES:
--
--    1.1.1.2 (3)
--
-- DESIGN UNIT ORDERING:
--
--    ENT00703(ARCH00703)
--    ENT00703_Test_Bench(ARCH00703_Test_Bench)
--
-- REVISION HISTORY:
--
--    25-JUN-1987   - initial revision
--
-- NOTES:
--
--    self-checking
--    automatically generated
--
use WORK.STANDARD_TYPES.all ;
entity ENT00703 is
   port (
          toggle : buffer switch ;
       i_st_rec1_1, i_st_rec1_2 : buffer st_rec1
          := c_st_rec1_1
          ;
       i_st_rec2_1, i_st_rec2_2 : buffer st_rec2
          := c_st_rec2_1
          ;
       i_st_rec3_1, i_st_rec3_2 : buffer st_rec3
          := c_st_rec3_1
          ;
       i_st_arr1_1, i_st_arr1_2 : buffer st_arr1
          := c_st_arr1_1
          ;
       i_st_arr2_1, i_st_arr2_2 : buffer st_arr2
          := c_st_arr2_1
          ;
       i_st_arr3_1, i_st_arr3_2 : buffer st_arr3
          := c_st_arr3_1
            ) ;
begin
end ENT00703 ;
--
architecture ARCH00703 of ENT00703 is
begin
   process
      variable correct : boolean := true ;
   begin
--
      toggle <= up ;
      i_st_rec1_1 <= c_st_rec1_2 ;
      i_st_rec1_2 <= c_st_rec1_2 ;
      i_st_rec2_1 <= c_st_rec2_2 ;
      i_st_rec2_2 <= c_st_rec2_2 ;
      i_st_rec3_1 <= c_st_rec3_2 ;
      i_st_rec3_2 <= c_st_rec3_2 ;
      i_st_arr1_1 <= c_st_arr1_2 ;
      i_st_arr1_2 <= c_st_arr1_2 ;
      i_st_arr2_1 <= c_st_arr2_2 ;
      i_st_arr2_2 <= c_st_arr2_2 ;
      i_st_arr3_1 <= c_st_arr3_2 ;
      i_st_arr3_2 <= c_st_arr3_2 ;
      test_report ( "ENT00703" ,
      "Open composite buffer ports with static subtypes" ,
      correct) ;
      wait ;
   end process ;
end ARCH00703 ;
--
use WORK.STANDARD_TYPES.all ;
entity ENT00703_Test_Bench is
end ENT00703_Test_Bench ;
--
architecture ARCH00703_Test_Bench of ENT00703_Test_Bench is
begin
   L1:
   block
--
      signal toggle : switch ;
--
      component UUT
      end component ;
--
      for CIS1 : UUT use entity WORK.ENT00703 ( ARCH00703 )
       port map (
                                       toggle ,
                               open, open,
                               open, open,
                               open, open,
                               open, open,
                               open, open,
                               open, open
                                      ) ;
--
   begin
      CIS1 : UUT ;
   end block L1 ;
end ARCH00703_Test_Bench ;
