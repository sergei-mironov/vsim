-------------------------------------------------------------------------------
	--
	--	   Copyright (c) 1989 by Intermetrics, Inc.
	--                All rights reserved.
	--
-------------------------------------------------------------------------------
--
-- TEST NAME:
--
--    CT00604
--
-- AUTHOR:
--
--    G. Tominovich
--
-- TEST OBJECTIVES:
--
--    11.1 (1)
--
-- DESIGN UNIT ORDERING:
--
--    N/A
--
-- REVISION HISTORY:
--
--    24-AUG-1987   - initial revision
--
-- NOTES:
--
--    will be used in conjunction with test ct00607
--
--
package body PKG00603 is
   procedure Proc is
   begin
      Null ;
   end Proc ;
end PKG00603 ;
--
